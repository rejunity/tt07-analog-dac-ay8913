magic
tech sky130A
magscale 1 2
timestamp 1716422392
<< metal1 >>
rect 21630 40950 21930 40956
rect 21630 40644 21930 40650
rect 30809 40800 31289 40806
rect 30809 40314 31289 40320
rect 20854 33800 20860 34400
rect 21460 33800 22260 34400
<< via1 >>
rect 21630 40650 21930 40950
rect 30809 40320 31289 40800
rect 20860 33800 21460 34400
<< metal2 >>
rect 20960 40954 23040 41000
rect 20955 40950 23040 40954
rect 20950 40945 21630 40950
rect 20950 40655 20955 40945
rect 21245 40655 21630 40945
rect 20950 40650 21630 40655
rect 21930 40650 23040 40950
rect 20955 40646 23040 40650
rect 20960 40600 23040 40646
rect 21151 40395 21813 40434
rect 21151 40233 21189 40395
rect 21351 40233 21813 40395
rect 30780 40320 30809 40800
rect 31289 40651 31460 40800
rect 31456 40484 31460 40651
rect 31289 40320 31460 40484
rect 21151 40195 21813 40233
rect 21151 39995 21815 40034
rect 21151 39833 21189 39995
rect 21351 39833 21815 39995
rect 21151 39795 21815 39833
rect 21151 39595 21807 39634
rect 21151 39433 21189 39595
rect 21351 39433 21807 39595
rect 21151 39395 21807 39433
rect 21151 39195 21815 39234
rect 21151 39033 21189 39195
rect 21351 39033 21815 39195
rect 21151 38995 21815 39033
rect 21151 38795 21813 38834
rect 21151 38633 21189 38795
rect 21351 38633 21813 38795
rect 21151 38595 21813 38633
rect 21151 38395 21819 38434
rect 21151 38233 21189 38395
rect 21351 38233 21819 38395
rect 21151 38195 21819 38233
rect 21151 37995 21821 38034
rect 21151 37833 21189 37995
rect 21351 37833 21821 37995
rect 21151 37795 21821 37833
rect 21151 37595 21819 37634
rect 21151 37433 21189 37595
rect 21351 37433 21819 37595
rect 21151 37395 21819 37433
rect 21151 37195 21815 37234
rect 21151 37033 21189 37195
rect 21351 37033 21815 37195
rect 21151 36995 21815 37033
rect 21151 36795 21815 36834
rect 21151 36633 21189 36795
rect 21351 36633 21815 36795
rect 21151 36595 21815 36633
rect 21151 36395 21817 36434
rect 21151 36233 21189 36395
rect 21351 36233 21817 36395
rect 21151 36195 21817 36233
rect 21151 35995 21811 36034
rect 21151 35833 21189 35995
rect 21351 35833 21811 35995
rect 21151 35795 21811 35833
rect 21149 35555 21815 35594
rect 21149 35393 21187 35555
rect 21349 35393 21815 35555
rect 21149 35355 21815 35393
rect 21151 35195 21817 35234
rect 21151 35033 21189 35195
rect 21351 35033 21817 35195
rect 21151 34995 21817 35033
rect 21151 34795 21815 34834
rect 21151 34633 21189 34795
rect 21351 34633 21815 34795
rect 21151 34595 21815 34633
rect 20860 34400 21460 34406
rect 20520 34245 20860 34400
rect 20520 33955 20555 34245
rect 20845 33955 20860 34245
rect 20520 33800 20860 33955
rect 20860 33794 21460 33800
<< via2 >>
rect 20955 40655 21245 40945
rect 21189 40233 21351 40395
rect 31289 40484 31456 40651
rect 21189 39833 21351 39995
rect 21189 39433 21351 39595
rect 21189 39033 21351 39195
rect 21189 38633 21351 38795
rect 21189 38233 21351 38395
rect 21189 37833 21351 37995
rect 21189 37433 21351 37595
rect 21189 37033 21351 37195
rect 21189 36633 21351 36795
rect 21189 36233 21351 36395
rect 21189 35833 21351 35995
rect 21187 35393 21349 35555
rect 21189 35033 21351 35195
rect 21189 34633 21351 34795
rect 20555 33955 20845 34245
<< metal3 >>
rect 17403 40950 17701 40955
rect 17402 40949 21250 40950
rect 17402 40651 17403 40949
rect 17701 40945 21250 40949
rect 17701 40655 20955 40945
rect 21245 40655 21250 40945
rect 31285 40656 31460 40661
rect 17701 40651 21250 40655
rect 17402 40650 21250 40651
rect 31284 40655 31461 40656
rect 17403 40645 17701 40650
rect 31284 40480 31285 40655
rect 31460 40480 31461 40655
rect 31284 40479 31461 40480
rect 31285 40474 31460 40479
rect 21076 40395 21356 40400
rect 21076 40346 21189 40395
rect 21076 40282 21130 40346
rect 21076 40233 21189 40282
rect 21351 40233 21356 40395
rect 21076 40228 21356 40233
rect 21076 39995 21356 40000
rect 21076 39946 21189 39995
rect 21076 39882 21130 39946
rect 21076 39833 21189 39882
rect 21351 39833 21356 39995
rect 21076 39828 21356 39833
rect 21076 39595 21356 39600
rect 21076 39546 21189 39595
rect 21076 39482 21130 39546
rect 21076 39433 21189 39482
rect 21351 39433 21356 39595
rect 21076 39428 21356 39433
rect 21076 39195 21356 39200
rect 21076 39146 21189 39195
rect 21076 39082 21130 39146
rect 21076 39033 21189 39082
rect 21351 39033 21356 39195
rect 21076 39028 21356 39033
rect 21076 38795 21356 38800
rect 21076 38746 21189 38795
rect 21076 38682 21130 38746
rect 21076 38633 21189 38682
rect 21351 38633 21356 38795
rect 21076 38628 21356 38633
rect 21076 38395 21356 38400
rect 21076 38346 21189 38395
rect 21076 38282 21130 38346
rect 21076 38233 21189 38282
rect 21351 38233 21356 38395
rect 21076 38228 21356 38233
rect 21076 37995 21356 38000
rect 21076 37946 21189 37995
rect 21076 37882 21130 37946
rect 21076 37833 21189 37882
rect 21351 37833 21356 37995
rect 21076 37828 21356 37833
rect 21076 37595 21356 37600
rect 21076 37546 21189 37595
rect 21076 37482 21130 37546
rect 21076 37433 21189 37482
rect 21351 37433 21356 37595
rect 21076 37428 21356 37433
rect 21076 37195 21356 37200
rect 21076 37146 21189 37195
rect 21076 37082 21130 37146
rect 21076 37033 21189 37082
rect 21351 37033 21356 37195
rect 21076 37028 21356 37033
rect 21076 36795 21356 36800
rect 21076 36746 21189 36795
rect 21076 36682 21130 36746
rect 21076 36633 21189 36682
rect 21351 36633 21356 36795
rect 21076 36628 21356 36633
rect 21076 36395 21356 36400
rect 21076 36346 21189 36395
rect 21076 36282 21130 36346
rect 21076 36233 21189 36282
rect 21351 36233 21356 36395
rect 21076 36228 21356 36233
rect 21076 35995 21356 36000
rect 21076 35946 21189 35995
rect 21076 35882 21130 35946
rect 21076 35833 21189 35882
rect 21351 35833 21356 35995
rect 21076 35828 21356 35833
rect 21074 35555 21354 35560
rect 21074 35506 21187 35555
rect 21074 35442 21128 35506
rect 21074 35393 21187 35442
rect 21349 35393 21354 35555
rect 21074 35388 21354 35393
rect 21076 35195 21356 35200
rect 21076 35146 21189 35195
rect 21076 35082 21130 35146
rect 21076 35033 21189 35082
rect 21351 35033 21356 35195
rect 21076 35028 21356 35033
rect 21076 34795 21356 34800
rect 21076 34746 21189 34795
rect 21076 34682 21130 34746
rect 21076 34633 21189 34682
rect 21351 34633 21356 34795
rect 21076 34628 21356 34633
rect 8951 34250 9249 34255
rect 8950 34249 20850 34250
rect 8950 33951 8951 34249
rect 9249 34245 20850 34249
rect 9249 33955 20555 34245
rect 20845 33955 20850 34245
rect 9249 33951 20850 33955
rect 8950 33950 20850 33951
rect 8951 33945 9249 33950
<< via3 >>
rect 17403 40651 17701 40949
rect 31285 40651 31460 40655
rect 31285 40484 31289 40651
rect 31289 40484 31456 40651
rect 31456 40484 31460 40651
rect 31285 40480 31460 40484
rect 21130 40282 21189 40346
rect 21189 40282 21194 40346
rect 21130 39882 21189 39946
rect 21189 39882 21194 39946
rect 21130 39482 21189 39546
rect 21189 39482 21194 39546
rect 21130 39082 21189 39146
rect 21189 39082 21194 39146
rect 21130 38682 21189 38746
rect 21189 38682 21194 38746
rect 21130 38282 21189 38346
rect 21189 38282 21194 38346
rect 21130 37882 21189 37946
rect 21189 37882 21194 37946
rect 21130 37482 21189 37546
rect 21189 37482 21194 37546
rect 21130 37082 21189 37146
rect 21189 37082 21194 37146
rect 21130 36682 21189 36746
rect 21189 36682 21194 36746
rect 21130 36282 21189 36346
rect 21189 36282 21194 36346
rect 21130 35882 21189 35946
rect 21189 35882 21194 35946
rect 21128 35442 21187 35506
rect 21187 35442 21192 35506
rect 21130 35082 21189 35146
rect 21189 35082 21194 35146
rect 21130 34682 21189 34746
rect 21189 34682 21194 34746
rect 8951 33951 9249 34249
<< metal4 >>
rect 798 44708 858 45152
rect 1534 44708 1594 45152
rect 2270 44708 2330 45152
rect 3006 44708 3066 45152
rect 3742 44708 3802 45152
rect 4478 44708 4538 45152
rect 5214 44708 5274 45152
rect 5950 44708 6010 45152
rect 6686 44708 6746 45152
rect 7422 44708 7482 45152
rect 8158 44708 8218 45152
rect 8894 44708 8954 45152
rect 9630 44708 9690 45152
rect 10366 44708 10426 45152
rect 11102 44708 11162 45152
rect 11838 44708 11898 45152
rect 12574 44708 12634 45152
rect 13310 44708 13370 45152
rect 14046 44708 14106 45152
rect 14782 44708 14842 45152
rect 15518 44708 15578 45152
rect 16254 44708 16314 45152
rect 16990 44708 17050 45152
rect 17726 44708 17786 45152
rect 798 44648 17786 44708
rect 200 34250 500 44152
rect 5950 44084 6010 44648
rect 9910 44152 9970 44648
rect 10366 44642 10426 44648
rect 9800 44084 10100 44152
rect 5950 44024 10100 44084
rect 9800 40950 10100 44024
rect 9800 40949 17702 40950
rect 9800 40651 17403 40949
rect 17701 40651 17702 40949
rect 9800 40650 17702 40651
rect 200 34249 9250 34250
rect 200 33951 8951 34249
rect 9249 33951 9250 34249
rect 200 33950 9250 33951
rect 200 1000 500 33950
rect 9800 1000 10100 40650
rect 18462 34744 18522 45152
rect 19198 43744 19258 45152
rect 18598 43720 19258 43744
rect 18598 43684 19256 43720
rect 18598 35144 18658 43684
rect 19934 43604 19994 45152
rect 18738 43544 19996 43604
rect 18738 35506 18798 43544
rect 19934 43542 19994 43544
rect 20670 43464 20730 45152
rect 18882 43404 20730 43464
rect 18882 35942 18942 43404
rect 20670 43402 20730 43404
rect 21406 43332 21466 45152
rect 19046 43272 21466 43332
rect 19046 36342 19106 43272
rect 22142 43210 22202 45152
rect 19206 43150 22202 43210
rect 19206 36742 19266 43150
rect 22878 43080 22938 45152
rect 19342 43020 22938 43080
rect 19342 37140 19402 43020
rect 23614 42956 23674 45152
rect 23014 42918 23674 42956
rect 19488 42858 23674 42918
rect 19488 37538 19548 42858
rect 24350 42792 24410 45152
rect 19628 42732 24410 42792
rect 19628 37940 19688 42732
rect 25086 42630 25146 45152
rect 19782 42570 25146 42630
rect 19782 38350 19842 42570
rect 25822 42438 25882 45152
rect 19920 42378 25882 42438
rect 19920 38742 19980 42378
rect 26558 42266 26618 45152
rect 20048 42206 26618 42266
rect 20048 39142 20108 42206
rect 27294 42096 27354 45152
rect 20186 42036 27354 42096
rect 20186 39544 20246 42036
rect 28030 41958 28090 45152
rect 20336 41898 28090 41958
rect 20336 39944 20396 41898
rect 28766 41808 28826 45152
rect 20474 41748 28826 41808
rect 20474 40334 20534 41748
rect 29502 41642 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 20618 41582 29562 41642
rect 20618 41312 20678 41582
rect 31284 40655 31461 40656
rect 31284 40480 31285 40655
rect 31460 40480 31461 40655
rect 21129 40346 21195 40347
rect 21129 40344 21130 40346
rect 20984 40334 21130 40344
rect 20474 40284 21130 40334
rect 20474 40274 21036 40284
rect 21129 40282 21130 40284
rect 21194 40282 21195 40346
rect 21129 40281 21195 40282
rect 21129 39946 21195 39947
rect 21129 39944 21130 39946
rect 20336 39884 21130 39944
rect 21129 39882 21130 39884
rect 21194 39882 21195 39946
rect 21129 39881 21195 39882
rect 21129 39546 21195 39547
rect 21129 39544 21130 39546
rect 20186 39484 21130 39544
rect 21129 39482 21130 39484
rect 21194 39482 21195 39546
rect 21129 39481 21195 39482
rect 21129 39146 21195 39147
rect 21129 39144 21130 39146
rect 20984 39142 21130 39144
rect 20048 39084 21130 39142
rect 20048 39082 21052 39084
rect 21129 39082 21130 39084
rect 21194 39082 21195 39146
rect 21129 39081 21195 39082
rect 21129 38746 21195 38747
rect 21129 38744 21130 38746
rect 20984 38742 21130 38744
rect 19920 38684 21130 38742
rect 19920 38682 21048 38684
rect 21129 38682 21130 38684
rect 21194 38682 21195 38746
rect 21129 38681 21195 38682
rect 19782 38344 21036 38350
rect 21129 38346 21195 38347
rect 21129 38344 21130 38346
rect 19782 38290 21130 38344
rect 20984 38284 21130 38290
rect 21129 38282 21130 38284
rect 21194 38282 21195 38346
rect 21129 38281 21195 38282
rect 21129 37946 21195 37947
rect 21129 37944 21130 37946
rect 20984 37940 21130 37944
rect 19628 37884 21130 37940
rect 19628 37880 21052 37884
rect 21129 37882 21130 37884
rect 21194 37882 21195 37946
rect 21129 37881 21195 37882
rect 21129 37546 21195 37547
rect 21129 37544 21130 37546
rect 20984 37538 21130 37544
rect 19488 37484 21130 37538
rect 19488 37478 21026 37484
rect 21129 37482 21130 37484
rect 21194 37482 21195 37546
rect 21129 37481 21195 37482
rect 21129 37146 21195 37147
rect 21129 37144 21130 37146
rect 20984 37140 21130 37144
rect 19342 37084 21130 37140
rect 19342 37080 21036 37084
rect 21129 37082 21130 37084
rect 21194 37082 21195 37146
rect 21129 37081 21195 37082
rect 21129 36746 21195 36747
rect 21129 36744 21130 36746
rect 20984 36742 21130 36744
rect 19206 36684 21130 36742
rect 19206 36682 21038 36684
rect 21129 36682 21130 36684
rect 21194 36682 21195 36746
rect 21129 36681 21195 36682
rect 21129 36346 21195 36347
rect 21129 36344 21130 36346
rect 20984 36342 21130 36344
rect 19046 36284 21130 36342
rect 19046 36282 21042 36284
rect 21129 36282 21130 36284
rect 21194 36282 21195 36346
rect 21129 36281 21195 36282
rect 21129 35946 21195 35947
rect 21129 35944 21130 35946
rect 20984 35942 21130 35944
rect 18882 35884 21130 35942
rect 18882 35882 21036 35884
rect 21129 35882 21130 35884
rect 21194 35882 21195 35946
rect 21129 35881 21195 35882
rect 21127 35506 21193 35507
rect 18738 35504 21060 35506
rect 21127 35504 21128 35506
rect 18738 35446 21128 35504
rect 20982 35444 21128 35446
rect 21127 35442 21128 35444
rect 21192 35442 21193 35506
rect 21127 35441 21193 35442
rect 21129 35146 21195 35147
rect 21129 35144 21130 35146
rect 18598 35084 21130 35144
rect 18598 35078 18658 35084
rect 21129 35082 21130 35084
rect 21194 35082 21195 35146
rect 21129 35081 21195 35082
rect 21129 34746 21195 34747
rect 21129 34744 21130 34746
rect 18462 34684 21130 34744
rect 21129 34682 21130 34684
rect 21194 34682 21195 34746
rect 21129 34681 21195 34682
rect 31284 200 31461 40480
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 200
use dac_16nfet  dac_16nfet_0
timestamp 1716419193
transform 1 0 21611 0 1 40600
box -11 -6800 9500 406
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31282 0 31462 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26866 0 27046 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22450 0 22630 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18034 0 18214 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13618 0 13798 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9202 0 9382 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4786 0 4966 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 370 0 550 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 4800 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 4800 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
