magic
tech sky130A
timestamp 1716300029
<< pwell >>
rect -173 -155 173 155
<< nmoslvt >>
rect -75 -50 75 50
<< ndiff >>
rect -104 44 -75 50
rect -104 -44 -98 44
rect -81 -44 -75 44
rect -104 -50 -75 -44
rect 75 44 104 50
rect 75 -44 81 44
rect 98 -44 104 44
rect 75 -50 104 -44
<< ndiffc >>
rect -98 -44 -81 44
rect 81 -44 98 44
<< psubdiff >>
rect -155 120 -107 137
rect 107 120 155 137
rect -155 89 -138 120
rect 138 89 155 120
rect -155 -120 -138 -89
rect 138 -120 155 -89
rect -155 -137 -107 -120
rect 107 -137 155 -120
<< psubdiffcont >>
rect -107 120 107 137
rect -155 -89 -138 89
rect 138 -89 155 89
rect -107 -137 107 -120
<< poly >>
rect -75 86 75 94
rect -75 69 -67 86
rect 67 69 75 86
rect -75 50 75 69
rect -75 -69 75 -50
rect -75 -86 -67 -69
rect 67 -86 75 -69
rect -75 -94 75 -86
<< polycont >>
rect -67 69 67 86
rect -67 -86 67 -69
<< locali >>
rect -155 120 -107 137
rect 107 120 155 137
rect -155 89 -138 120
rect 138 89 155 120
rect -75 69 -67 86
rect 67 69 75 86
rect -98 44 -81 52
rect -98 -52 -81 -44
rect 81 44 98 52
rect 81 -52 98 -44
rect -75 -86 -67 -69
rect 67 -86 75 -69
rect -155 -120 -138 -89
rect 138 -120 155 -89
rect -155 -137 -107 -120
rect 107 -137 155 -120
<< viali >>
rect -67 69 67 86
rect -98 -44 -81 44
rect 81 -44 98 44
rect -67 -86 67 -69
<< metal1 >>
rect -73 86 73 89
rect -73 69 -67 86
rect 67 69 73 86
rect -73 66 73 69
rect -101 44 -78 50
rect -101 -44 -98 44
rect -81 -44 -78 44
rect -101 -50 -78 -44
rect 78 44 101 50
rect 78 -44 81 44
rect 98 -44 101 44
rect 78 -50 101 -44
rect -73 -69 73 -66
rect -73 -86 -67 -69
rect 67 -86 73 -69
rect -73 -89 73 -86
<< properties >>
string FIXED_BBOX -146 -128 146 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 1.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
