magic
tech sky130A
magscale 1 2
timestamp 1716419193
<< pwell >>
rect 3980 -200 4100 -140
rect 2370 -2340 2660 -2000
rect 4820 -3616 5050 -3614
rect 5536 -3616 5766 -3614
rect 6252 -3616 6482 -3614
rect 6968 -3616 7198 -3614
rect 7684 -3616 7914 -3614
rect 4812 -3618 5060 -3616
rect 5528 -3618 5776 -3616
rect 6244 -3618 6492 -3616
rect 6960 -3618 7208 -3616
rect 7676 -3618 7924 -3616
rect 4806 -4228 5060 -3618
rect 5522 -4228 5776 -3618
rect 6238 -4228 6492 -3618
rect 6954 -4228 7208 -3618
rect 7670 -4228 7924 -3618
<< locali >>
rect 532 -178 640 -144
rect 1000 -178 3088 -144
<< viali >>
rect 640 -180 1000 -140
rect 3560 -580 3920 -540
rect 5760 -880 6140 -840
rect 7400 -1280 7760 -1240
rect 2340 -2070 2650 -2030
rect 2420 -2320 2650 -2280
rect 3170 -2920 3380 -2880
rect 3070 -3540 3380 -3500
rect 4380 -3590 4470 -3540
rect 3070 -3660 3380 -3620
rect 3860 -3650 4080 -3610
rect 4290 -3710 4340 -3630
rect 4820 -4188 4854 -3636
rect 5016 -4196 5050 -3644
rect 5536 -4188 5570 -3636
rect 5732 -4196 5766 -3644
rect 6252 -4188 6286 -3636
rect 6448 -4196 6482 -3644
rect 6968 -4188 7002 -3636
rect 7164 -4196 7198 -3644
rect 7684 -4188 7718 -3636
rect 7880 -4196 7914 -3644
rect 8390 -6170 8430 -5620
<< metal1 >>
rect 620 400 1020 406
rect 0 0 620 400
rect 620 -140 1020 0
rect 620 -180 640 -140
rect 1000 -180 1020 -140
rect 620 -200 1020 -180
rect 1080 -100 9500 200
rect 1080 -160 5100 -100
rect 1080 -200 3480 -160
rect 0 -320 200 -200
rect 1080 -237 3000 -200
rect 622 -292 3000 -237
rect -3 -490 3 -320
rect 173 -400 200 -320
rect 407 -320 577 -314
rect 173 -490 179 -400
rect 407 -496 577 -490
rect 3047 -320 3217 -314
rect 3047 -496 3217 -490
rect 2412 -516 2998 -510
rect 0 -720 200 -600
rect 168 -800 200 -720
rect 0 -894 168 -888
rect 622 -900 2998 -516
rect 3534 -600 3540 -200
rect 3940 -600 3946 -200
rect 4020 -300 5100 -160
rect 5300 -300 9500 -100
rect 4020 -400 9500 -300
rect 4020 -520 5680 -400
rect 4020 -640 5192 -520
rect 3522 -692 5192 -640
rect 3620 -698 3980 -692
rect 3306 -720 3474 -714
rect 3306 -894 3474 -888
rect 5232 -720 5400 -714
rect 5232 -894 5400 -888
rect 5734 -900 5740 -500
rect 6140 -900 6146 -500
rect 6200 -600 6800 -400
rect 0 -1022 200 -1000
rect 0 -1186 4 -1022
rect 168 -1186 200 -1022
rect 0 -1200 200 -1186
rect 600 -1096 2998 -900
rect -11 -1499 -5 -1337
rect 157 -1400 163 -1337
rect 157 -1499 200 -1400
rect 0 -1600 200 -1499
rect -1 -1880 5 -1730
rect 155 -1800 161 -1730
rect 155 -1880 200 -1800
rect 0 -2000 200 -1880
rect 0 -2259 200 -2200
rect -5 -2265 200 -2259
rect 145 -2400 200 -2265
rect -5 -2421 145 -2415
rect 0 -2710 200 -2600
rect 0 -2800 15 -2710
rect 165 -2800 200 -2710
rect 15 -2866 165 -2860
rect 600 -2850 1200 -1096
rect 2412 -1120 2998 -1096
rect 3522 -916 3882 -910
rect 3522 -1120 5192 -916
rect 6200 -940 6892 -600
rect 7000 -780 9500 -400
rect 7840 -842 8240 -780
rect 5726 -992 6892 -940
rect 2412 -1270 5192 -1120
rect 5522 -1022 5686 -1016
rect 5522 -1192 5686 -1186
rect 6948 -1022 7112 -1016
rect 6948 -1192 7112 -1186
rect 2412 -1320 5180 -1270
rect 5726 -1320 6892 -1212
rect 7374 -1300 7380 -900
rect 7780 -1300 7786 -900
rect 2412 -1480 6892 -1320
rect 7840 -1340 8242 -842
rect 7426 -1390 8242 -1340
rect 2412 -1693 2998 -1480
rect 4820 -1632 6892 -1480
rect 7211 -1424 7373 -1418
rect 7211 -1592 7373 -1586
rect 8291 -1424 8453 -1418
rect 8291 -1592 8453 -1586
rect 7426 -1614 7978 -1610
rect 4820 -1680 6880 -1632
rect 2225 -1730 2375 -1724
rect 2225 -1886 2375 -1880
rect 3055 -1730 3205 -1724
rect 3055 -1886 3205 -1880
rect 5924 -1762 6776 -1680
rect 7426 -1762 8242 -1614
rect 2700 -1990 3000 -1920
rect 2320 -2030 2670 -2000
rect 2320 -2070 2340 -2030
rect 2650 -2070 2670 -2030
rect 2320 -2310 2350 -2070
rect 2630 -2280 2670 -2070
rect 2320 -2320 2420 -2310
rect 2650 -2320 2670 -2280
rect 2320 -2340 2670 -2320
rect 2700 -2240 5730 -1990
rect 5924 -2160 8242 -1762
rect 8520 -2240 9500 -780
rect 2700 -2260 9500 -2240
rect 2700 -2430 2910 -2260
rect 2946 -2264 9500 -2260
rect 3180 -2440 3400 -2430
rect 2416 -2480 2545 -2474
rect 2875 -2480 3004 -2474
rect 2410 -2609 2416 -2480
rect 2545 -2609 2551 -2480
rect 2416 -2615 2545 -2609
rect 2875 -2615 3004 -2609
rect 3174 -2660 3180 -2440
rect 3400 -2660 3406 -2440
rect 2510 -2850 2910 -2660
rect 0 -3140 200 -3000
rect 0 -3200 15 -3140
rect 165 -3200 200 -3140
rect 600 -3080 2910 -2850
rect 3150 -2880 3400 -2660
rect 3150 -2920 3170 -2880
rect 3380 -2920 3400 -2880
rect 3150 -2930 3400 -2920
rect 15 -3296 165 -3290
rect 600 -3250 3110 -3080
rect 3150 -3104 3156 -2976
rect 3284 -3104 3290 -2976
rect 4150 -3080 9500 -2264
rect 0 -3510 200 -3400
rect 0 -3600 5 -3510
rect 155 -3600 200 -3510
rect 5 -3666 155 -3660
rect 0 -3875 200 -3800
rect -1 -4025 5 -3875
rect 155 -4000 200 -3875
rect 155 -4025 161 -4000
rect 0 -4285 200 -4200
rect 0 -4400 5 -4285
rect 155 -4400 200 -4285
rect 5 -4441 155 -4435
rect 0 -4675 200 -4600
rect -11 -4825 -5 -4675
rect 145 -4800 200 -4675
rect 145 -4825 151 -4800
rect 0 -5048 200 -5000
rect -5 -5054 200 -5048
rect 145 -5200 200 -5054
rect -5 -5210 145 -5204
rect 0 -5485 200 -5400
rect 0 -5600 15 -5485
rect 9 -5635 15 -5600
rect 165 -5600 200 -5485
rect 165 -5635 171 -5600
rect 0 -5835 200 -5800
rect -11 -5985 -5 -5835
rect 145 -5985 200 -5835
rect 0 -6000 200 -5985
rect 600 -6200 1200 -3250
rect 2510 -3340 3110 -3250
rect 3156 -3326 3284 -3104
rect 2510 -3820 2910 -3340
rect 3150 -3454 3156 -3326
rect 3284 -3454 3290 -3326
rect 3340 -3338 9500 -3080
rect 3340 -3340 8504 -3338
rect 3050 -3500 3400 -3490
rect 3050 -3540 3070 -3500
rect 3380 -3540 3400 -3500
rect 3050 -3620 3400 -3540
rect 3050 -3660 3070 -3620
rect 3380 -3660 3400 -3620
rect 3050 -3670 3400 -3660
rect 2510 -3980 3110 -3820
rect 3159 -3846 3165 -3715
rect 3296 -3846 3302 -3715
rect 3440 -3820 3595 -3340
rect 3854 -3580 3860 -3370
rect 3850 -3590 3860 -3580
rect 4080 -3400 4086 -3370
rect 4080 -3540 4490 -3400
rect 4080 -3590 4380 -3540
rect 4470 -3590 4490 -3540
rect 3850 -3600 4490 -3590
rect 3850 -3610 4090 -3600
rect 3850 -3650 3860 -3610
rect 4080 -3650 4090 -3610
rect 3850 -3670 4090 -3650
rect 4270 -3630 4360 -3600
rect 4270 -3710 4290 -3630
rect 4340 -3710 4360 -3630
rect 4520 -3660 4680 -3340
rect 4820 -3616 5050 -3614
rect 4812 -3618 5060 -3616
rect 4480 -3710 4680 -3660
rect 4806 -3636 5060 -3618
rect 3835 -3725 3985 -3719
rect 4270 -3720 4360 -3710
rect 3159 -4085 3165 -3954
rect 3296 -4085 3302 -3954
rect 3340 -3990 3740 -3820
rect 4615 -3755 4762 -3749
rect 3835 -3881 3985 -3875
rect 3779 -4105 3785 -3955
rect 3935 -4105 3941 -3955
rect 4030 -4000 4250 -3800
rect 4289 -3905 4295 -3755
rect 4040 -4010 4250 -4000
rect 4070 -4358 4250 -4010
rect 4295 -3945 4370 -3905
rect 4295 -4100 4370 -4075
rect 4445 -4100 4451 -3755
rect 4615 -4100 4762 -4084
rect 4295 -4121 4451 -4100
rect 4068 -6200 4268 -4358
rect 4480 -6200 4680 -4169
rect 4806 -4188 4820 -3636
rect 4854 -3644 5060 -3636
rect 4854 -3729 5016 -3644
rect 4854 -3879 4860 -3729
rect 5010 -3879 5016 -3729
rect 4854 -4188 5016 -3879
rect 4806 -4196 5016 -4188
rect 5050 -4196 5060 -3644
rect 5184 -3722 5392 -3340
rect 5640 -3344 6106 -3340
rect 5536 -3616 5766 -3614
rect 5528 -3618 5776 -3616
rect 5522 -3636 5776 -3618
rect 5323 -3779 5473 -3773
rect 5097 -3929 5103 -3779
rect 5253 -3929 5259 -3779
rect 5323 -3935 5473 -3929
rect 4806 -4228 5060 -4196
rect 5522 -4188 5536 -3636
rect 5570 -3644 5776 -3636
rect 5570 -3729 5732 -3644
rect 5570 -3879 5576 -3729
rect 5726 -3879 5732 -3729
rect 5570 -4188 5732 -3879
rect 5522 -4196 5732 -4188
rect 5766 -4196 5776 -3644
rect 5906 -3716 6106 -3344
rect 6252 -3616 6482 -3614
rect 6244 -3618 6492 -3616
rect 6238 -3636 6492 -3618
rect 6045 -3767 6195 -3761
rect 5818 -3917 5824 -3767
rect 5974 -3917 5980 -3767
rect 6045 -3923 6195 -3917
rect 5522 -4228 5776 -4196
rect 6238 -4188 6252 -3636
rect 6286 -3644 6492 -3636
rect 6286 -3729 6448 -3644
rect 6286 -3879 6292 -3729
rect 6442 -3879 6448 -3729
rect 6286 -4188 6448 -3879
rect 6238 -4196 6448 -4188
rect 6482 -4196 6492 -3644
rect 6620 -3690 6820 -3340
rect 6968 -3616 7198 -3614
rect 6960 -3618 7208 -3616
rect 6954 -3636 7208 -3618
rect 6761 -3741 6911 -3735
rect 6530 -3891 6536 -3741
rect 6686 -3891 6692 -3741
rect 6761 -3897 6911 -3891
rect 6238 -4228 6492 -4196
rect 6954 -4188 6968 -3636
rect 7002 -3644 7208 -3636
rect 7002 -3729 7164 -3644
rect 7002 -3879 7008 -3729
rect 7158 -3879 7164 -3729
rect 7002 -4188 7164 -3879
rect 6954 -4196 7164 -4188
rect 7198 -4196 7208 -3644
rect 7340 -3692 7540 -3340
rect 7684 -3616 7914 -3614
rect 7676 -3618 7924 -3616
rect 7670 -3636 7924 -3618
rect 7475 -3737 7625 -3731
rect 7242 -3887 7248 -3737
rect 7398 -3887 7404 -3737
rect 7475 -3893 7625 -3887
rect 6954 -4228 7208 -4196
rect 7670 -4188 7684 -3636
rect 7718 -3644 7924 -3636
rect 7718 -3729 7880 -3644
rect 7718 -3879 7724 -3729
rect 7874 -3879 7880 -3729
rect 7718 -4188 7880 -3879
rect 7670 -4196 7880 -4188
rect 7914 -4196 7924 -3644
rect 8052 -3698 8252 -3340
rect 8195 -3743 8345 -3737
rect 7962 -3893 7968 -3743
rect 8118 -3893 8124 -3743
rect 8195 -3899 8345 -3893
rect 7670 -4228 7924 -4196
rect 5190 -6200 5392 -4350
rect 5819 -4537 5825 -4387
rect 5975 -4537 5981 -4387
rect 6039 -4553 6045 -4403
rect 6195 -4553 6201 -4403
rect 5908 -6200 6094 -4582
rect 6537 -4715 6687 -4709
rect 6755 -4865 6761 -4715
rect 6911 -4865 6917 -4715
rect 6537 -4871 6687 -4865
rect 6624 -6200 6810 -4904
rect 7251 -5221 7401 -5215
rect 7469 -5371 7475 -5221
rect 7625 -5371 7631 -5221
rect 7251 -5377 7401 -5371
rect 7340 -6200 7526 -5416
rect 8380 -5620 8710 -5600
rect 7969 -5925 8119 -5919
rect 8189 -6075 8195 -5925
rect 8345 -6075 8351 -5925
rect 7969 -6081 8119 -6075
rect -10 -6344 7800 -6200
rect 8056 -6344 8252 -6118
rect 8380 -6170 8390 -5620
rect 8430 -5890 8710 -5620
rect 8380 -6230 8710 -6170
rect 8430 -6260 8710 -6230
rect -10 -6548 8252 -6344
rect -10 -6800 7800 -6548
<< via1 >>
rect 620 0 1020 400
rect 3 -490 173 -320
rect 407 -490 577 -320
rect 3047 -490 3217 -320
rect 0 -888 168 -720
rect 3540 -540 3940 -200
rect 3540 -580 3560 -540
rect 3560 -580 3920 -540
rect 3920 -580 3940 -540
rect 3540 -600 3940 -580
rect 3306 -888 3474 -720
rect 5232 -888 5400 -720
rect 5740 -840 6140 -500
rect 5740 -880 5760 -840
rect 5760 -880 6140 -840
rect 5740 -900 6140 -880
rect 4 -1186 168 -1022
rect -5 -1499 157 -1337
rect 5 -1880 155 -1730
rect -5 -2415 145 -2265
rect 15 -2860 165 -2710
rect 5522 -1186 5686 -1022
rect 6948 -1186 7112 -1022
rect 7380 -1240 7780 -900
rect 7380 -1280 7400 -1240
rect 7400 -1280 7760 -1240
rect 7760 -1280 7780 -1240
rect 7380 -1300 7780 -1280
rect 7211 -1586 7373 -1424
rect 8291 -1586 8453 -1424
rect 2225 -1880 2375 -1730
rect 3055 -1880 3205 -1730
rect 2350 -2070 2630 -2030
rect 2350 -2280 2630 -2070
rect 2350 -2310 2420 -2280
rect 2420 -2310 2630 -2280
rect 2416 -2609 2545 -2480
rect 2875 -2609 3004 -2480
rect 3180 -2660 3400 -2440
rect 15 -3290 165 -3140
rect 3156 -3104 3284 -2976
rect 5 -3660 155 -3510
rect 5 -4025 155 -3875
rect 5 -4435 155 -4285
rect -5 -4825 145 -4675
rect -5 -5204 145 -5054
rect 15 -5635 165 -5485
rect -5 -5985 145 -5835
rect 3156 -3454 3284 -3326
rect 3165 -3846 3296 -3715
rect 3860 -3590 4080 -3370
rect 3165 -4085 3296 -3954
rect 3835 -3875 3985 -3725
rect 3785 -4105 3935 -3955
rect 4295 -3905 4445 -3755
rect 4370 -3945 4445 -3905
rect 4295 -4075 4445 -3945
rect 4370 -4100 4445 -4075
rect 4615 -4084 4762 -3755
rect 4860 -3879 5010 -3729
rect 5103 -3929 5253 -3779
rect 5323 -3929 5473 -3779
rect 5576 -3879 5726 -3729
rect 5824 -3917 5974 -3767
rect 6045 -3917 6195 -3767
rect 6292 -3879 6442 -3729
rect 6536 -3891 6686 -3741
rect 6761 -3891 6911 -3741
rect 7008 -3879 7158 -3729
rect 7248 -3887 7398 -3737
rect 7475 -3887 7625 -3737
rect 7724 -3879 7874 -3729
rect 7968 -3893 8118 -3743
rect 8195 -3893 8345 -3743
rect 5825 -4537 5975 -4387
rect 6045 -4553 6195 -4403
rect 6537 -4865 6687 -4715
rect 6761 -4865 6911 -4715
rect 7251 -5371 7401 -5221
rect 7475 -5371 7625 -5221
rect 7969 -6075 8119 -5925
rect 8195 -6075 8345 -5925
rect 8430 -6170 8710 -5890
<< metal2 >>
rect 600 0 620 400
rect 1020 0 8942 400
rect 3540 -200 3940 0
rect 3 -320 173 -314
rect 173 -490 407 -320
rect 577 -490 3047 -320
rect 3217 -490 3311 -320
rect 3 -496 173 -490
rect 3540 -606 3940 -600
rect 5740 -500 6140 0
rect -6 -888 0 -720
rect 168 -888 3306 -720
rect 3474 -888 5232 -720
rect 5400 -888 5407 -720
rect 5740 -906 6140 -900
rect 7380 -900 7780 0
rect -2 -1186 4 -1022
rect 168 -1186 5522 -1022
rect 5686 -1186 6948 -1022
rect 7112 -1186 7136 -1022
rect 7380 -1306 7780 -1300
rect -5 -1337 157 -1331
rect 157 -1424 3597 -1337
rect 157 -1499 7211 -1424
rect -5 -1505 157 -1499
rect 3435 -1586 7211 -1499
rect 7373 -1586 8291 -1424
rect 8453 -1586 8485 -1424
rect 5 -1730 155 -1724
rect 155 -1880 2225 -1730
rect 2375 -1880 3055 -1730
rect 3205 -1880 3211 -1730
rect 5 -1886 155 -1880
rect 8542 -2030 8942 0
rect -11 -2415 -5 -2265
rect 145 -2415 545 -2265
rect 2344 -2310 2350 -2030
rect 2630 -2310 8942 -2030
rect 395 -2470 545 -2415
rect 3180 -2440 3400 -2310
rect 395 -2480 3035 -2470
rect 395 -2609 2416 -2480
rect 2545 -2609 2875 -2480
rect 3004 -2609 3035 -2480
rect 395 -2620 3035 -2609
rect 3180 -2666 3400 -2660
rect 0 -2860 15 -2710
rect 165 -2860 3285 -2710
rect 3156 -2976 3284 -2860
rect 0 -3290 15 -3140
rect 165 -3290 2475 -3140
rect -1 -3660 5 -3510
rect 155 -3660 2175 -3510
rect 5 -3870 155 -3869
rect 0 -3875 155 -3870
rect 0 -4025 5 -3875
rect 155 -4025 1865 -3985
rect 0 -4135 1865 -4025
rect -1 -4435 5 -4285
rect 155 -4435 1525 -4285
rect 1375 -4550 1525 -4435
rect 1715 -4355 1865 -4135
rect 2025 -4145 2175 -3660
rect 2325 -3565 2475 -3290
rect 3156 -3326 3284 -3104
rect 3156 -3460 3284 -3454
rect 3860 -3064 4080 -2310
rect 8540 -3064 8942 -2310
rect 3860 -3344 8942 -3064
rect 3860 -3370 4080 -3344
rect 2325 -3715 3305 -3565
rect 3860 -3596 4080 -3590
rect 2325 -3720 2475 -3715
rect 3165 -3954 3296 -3846
rect 3165 -4091 3296 -4085
rect 3745 -3875 3835 -3725
rect 3985 -3875 3995 -3725
rect 4860 -3729 5010 -3344
rect 3745 -3955 3995 -3875
rect 4295 -3755 4762 -3735
rect 4295 -3945 4370 -3905
rect 3745 -4105 3785 -3955
rect 3935 -4105 3995 -3955
rect 4289 -4075 4295 -3945
rect 3745 -4145 3995 -4105
rect 2025 -4295 3995 -4145
rect 4295 -4100 4370 -4075
rect 4445 -4084 4615 -3755
rect 5576 -3729 5726 -3344
rect 4860 -3885 5010 -3879
rect 5100 -3779 5477 -3751
rect 4445 -4090 4762 -4084
rect 5100 -3929 5103 -3779
rect 5253 -3929 5323 -3779
rect 5473 -3929 5479 -3779
rect 6292 -3729 6442 -3344
rect 5576 -3885 5726 -3879
rect 5824 -3767 5974 -3751
rect 5974 -3917 6045 -3767
rect 6195 -3917 6201 -3767
rect 7008 -3729 7158 -3344
rect 6292 -3885 6442 -3879
rect 6536 -3741 6686 -3735
rect 6686 -3891 6761 -3741
rect 6911 -3891 6917 -3741
rect 7724 -3729 7874 -3344
rect 7008 -3885 7158 -3879
rect 7248 -3737 7398 -3731
rect 7398 -3887 7475 -3737
rect 7625 -3887 7631 -3737
rect 7724 -3885 7874 -3879
rect 7968 -3743 8118 -3737
rect 4445 -4100 4615 -4090
rect 4295 -4355 4445 -4100
rect 1715 -4505 4445 -4355
rect 5100 -4157 5253 -3929
rect 5327 -4157 5477 -3929
rect 5100 -4307 5477 -4157
rect 5824 -4087 5974 -3917
rect 5100 -4550 5250 -4307
rect 5824 -4387 5975 -4087
rect 5824 -4537 5825 -4387
rect 6045 -4403 6195 -3917
rect 5975 -4537 6045 -4403
rect -5 -4675 145 -4669
rect 1375 -4700 5255 -4550
rect 5824 -4553 6045 -4537
rect 5824 -4802 5974 -4553
rect 6045 -4559 6195 -4553
rect 6536 -4715 6686 -3891
rect 6761 -4715 6911 -3891
rect 145 -4825 5974 -4802
rect -5 -4952 5974 -4825
rect 6531 -4865 6537 -4715
rect 6687 -4865 6761 -4715
rect 6536 -5054 6686 -4865
rect 6761 -4871 6911 -4865
rect -11 -5204 -5 -5054
rect 145 -5204 6686 -5054
rect 7248 -5221 7398 -3887
rect 7475 -5221 7625 -3887
rect 7245 -5371 7251 -5221
rect 7401 -5371 7475 -5221
rect 15 -5485 165 -5479
rect 7248 -5570 7398 -5371
rect 7475 -5377 7625 -5371
rect 8118 -3893 8195 -3743
rect 8345 -3893 8351 -3743
rect 165 -5635 7398 -5570
rect 15 -5720 7398 -5635
rect -5 -5835 145 -5829
rect 7968 -5925 8118 -3893
rect 8195 -5925 8345 -3893
rect 8542 -5890 8942 -3344
rect -5 -6175 145 -5985
rect 7963 -6075 7969 -5925
rect 8119 -6075 8195 -5925
rect 7968 -6175 8118 -6075
rect 8195 -6081 8345 -6075
rect 8424 -6170 8430 -5890
rect 8710 -6170 8942 -5890
rect -5 -6325 8118 -6175
rect 8542 -6180 8942 -6170
rect 7968 -6342 8118 -6325
use sky130_fd_pr__nfet_01v8_lvt_PXK84T  XM1
timestamp 1716300029
transform 0 -1 8154 1 0 -4908
box -1396 -310 1396 310
use sky130_fd_pr__nfet_01v8_lvt_DV472Z  XM2
timestamp 1716300029
transform 0 -1 7438 1 0 -4554
box -1044 -310 1044 310
use sky130_fd_pr__nfet_01v8_lvt_S4XANK  XM3
timestamp 1716300029
transform 0 -1 6722 1 0 -4302
box -796 -310 796 310
use sky130_fd_pr__nfet_01v8_lvt_XA7BLB  XM4
timestamp 1716300029
transform 0 1 1810 -1 0 -404
box -296 -1410 296 1410
use sky130_fd_pr__nfet_01v8_lvt_PVCJZS  XM5
timestamp 1716300029
transform 0 -1 6006 1 0 -4152
box -620 -310 620 310
use sky130_fd_pr__nfet_01v8_lvt_V433WY  XM6
timestamp 1716300029
transform 0 -1 5290 1 0 -4034
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_lvt_NWFTZM  XM7
timestamp 1716300029
transform 0 1 4580 1 0 -3912
box -408 -310 408 310
use sky130_fd_pr__nfet_01v8_lvt_UJ7Z4X  XM8
timestamp 1716300029
transform -1 0 3226 0 -1 -3210
box -296 -360 296 360
use sky130_fd_pr__nfet_01v8_lvt_C8TQ3N  XM9
timestamp 1716300029
transform 0 1 2710 -1 0 -1804
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_lvt_XESRVR  XM10
timestamp 1716300029
transform 0 1 2712 -1 0 -2544
box -296 -422 296 422
use sky130_fd_pr__nfet_01v8_lvt_N5KR3K  XM11
timestamp 1716300029
transform 1 0 3866 0 1 -3900
box -346 -310 346 310
use sky130_fd_pr__nfet_01v8_lvt_69TQ3K  XM12
timestamp 1716300029
transform 1 0 3226 0 1 -3900
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_lvt_P5KZ23  XM14
timestamp 1716300029
transform 0 1 4358 -1 0 -804
box -296 -1058 296 1058
use sky130_fd_pr__nfet_01v8_lvt_HQ7AL5  XM15
timestamp 1716300029
transform 0 1 6310 -1 0 -1104
box -296 -810 296 810
use sky130_fd_pr__nfet_01v8_lvt_L27GYG  XM16
timestamp 1716300029
transform 0 1 7834 -1 0 -1504
box -296 -634 296 634
<< labels >>
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 AT0
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 AT1
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 AT2
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 AT3
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 AT4
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 AT5
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 AT6
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 AT7
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 AT8
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 AT9
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 AT10
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 AT11
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 AT12
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 AT13
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 AT14
port 15 nsew
flabel metal1 9300 0 9500 200 0 FreeSans 256 0 0 0 OUT
port 16 nsew
flabel metal1 20 180 220 380 0 FreeSans 256 0 0 0 VSS
port 17 nsew
flabel metal1 600 -6800 800 -6600 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
