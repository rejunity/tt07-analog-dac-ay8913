magic
tech sky130A
timestamp 1716300029
<< pwell >>
rect -148 -211 148 211
<< nmoslvt >>
rect -50 -106 50 106
<< ndiff >>
rect -79 100 -50 106
rect -79 -100 -73 100
rect -56 -100 -50 100
rect -79 -106 -50 -100
rect 50 100 79 106
rect 50 -100 56 100
rect 73 -100 79 100
rect 50 -106 79 -100
<< ndiffc >>
rect -73 -100 -56 100
rect 56 -100 73 100
<< psubdiff >>
rect -130 176 -82 193
rect 82 176 130 193
rect -130 145 -113 176
rect 113 145 130 176
rect -130 -176 -113 -145
rect 113 -176 130 -145
rect -130 -193 -82 -176
rect 82 -193 130 -176
<< psubdiffcont >>
rect -82 176 82 193
rect -130 -145 -113 145
rect 113 -145 130 145
rect -82 -193 82 -176
<< poly >>
rect -50 142 50 150
rect -50 125 -42 142
rect 42 125 50 142
rect -50 106 50 125
rect -50 -125 50 -106
rect -50 -142 -42 -125
rect 42 -142 50 -125
rect -50 -150 50 -142
<< polycont >>
rect -42 125 42 142
rect -42 -142 42 -125
<< locali >>
rect -130 176 -82 193
rect 82 176 130 193
rect -130 145 -113 176
rect 113 145 130 176
rect -50 125 -42 142
rect 42 125 50 142
rect -73 100 -56 108
rect -73 -108 -56 -100
rect 56 100 73 108
rect 56 -108 73 -100
rect -50 -142 -42 -125
rect 42 -142 50 -125
rect -130 -176 -113 -145
rect 113 -176 130 -145
rect -130 -193 -82 -176
rect 82 -193 130 -176
<< viali >>
rect -42 125 42 142
rect -73 -100 -56 100
rect 56 -100 73 100
rect -42 -142 42 -125
<< metal1 >>
rect -48 142 48 145
rect -48 125 -42 142
rect 42 125 48 142
rect -48 122 48 125
rect -76 100 -53 106
rect -76 -100 -73 100
rect -56 -100 -53 100
rect -76 -106 -53 -100
rect 53 100 76 106
rect 53 -100 56 100
rect 73 -100 76 100
rect 53 -106 76 -100
rect -48 -125 48 -122
rect -48 -142 -42 -125
rect 42 -142 48 -125
rect -48 -145 48 -142
<< properties >>
string FIXED_BBOX -121 -184 121 184
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.12 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
