magic
tech sky130A
timestamp 1716300029
<< pwell >>
rect -698 -155 698 155
<< nmoslvt >>
rect -600 -50 600 50
<< ndiff >>
rect -629 44 -600 50
rect -629 -44 -623 44
rect -606 -44 -600 44
rect -629 -50 -600 -44
rect 600 44 629 50
rect 600 -44 606 44
rect 623 -44 629 44
rect 600 -50 629 -44
<< ndiffc >>
rect -623 -44 -606 44
rect 606 -44 623 44
<< psubdiff >>
rect -680 120 -632 137
rect 632 120 680 137
rect -680 89 -663 120
rect 663 89 680 120
rect -680 -120 -663 -89
rect 663 -120 680 -89
rect -680 -137 -632 -120
rect 632 -137 680 -120
<< psubdiffcont >>
rect -632 120 632 137
rect -680 -89 -663 89
rect 663 -89 680 89
rect -632 -137 632 -120
<< poly >>
rect -600 86 600 94
rect -600 69 -592 86
rect 592 69 600 86
rect -600 50 600 69
rect -600 -69 600 -50
rect -600 -86 -592 -69
rect 592 -86 600 -69
rect -600 -94 600 -86
<< polycont >>
rect -592 69 592 86
rect -592 -86 592 -69
<< locali >>
rect -680 120 -632 137
rect 632 120 680 137
rect -680 89 -663 120
rect 663 89 680 120
rect -600 69 -592 86
rect 592 69 600 86
rect -623 44 -606 52
rect -623 -52 -606 -44
rect 606 44 623 52
rect 606 -52 623 -44
rect -600 -86 -592 -69
rect 592 -86 600 -69
rect -680 -120 -663 -89
rect 663 -120 680 -89
rect -680 -137 -632 -120
rect 632 -137 680 -120
<< viali >>
rect -592 69 592 86
rect -623 -44 -606 44
rect 606 -44 623 44
rect -592 -86 592 -69
<< metal1 >>
rect -598 86 598 89
rect -598 69 -592 86
rect 592 69 598 86
rect -598 66 598 69
rect -626 44 -603 50
rect -626 -44 -623 44
rect -606 -44 -603 44
rect -626 -50 -603 -44
rect 603 44 626 50
rect 603 -44 606 44
rect 623 -44 626 44
rect 603 -50 626 -44
rect -598 -69 598 -66
rect -598 -86 -592 -69
rect 592 -86 598 -69
rect -598 -89 598 -86
<< properties >>
string FIXED_BBOX -671 -128 671 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 12.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
