MACRO tt_um_rejunity_analog_dac_ay8913
  CLASS BLOCK ;
  FOREIGN tt_um_rejunity_analog_dac_ay8913 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.148600 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.480000 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.240000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.120000 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.000000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.120000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.000000 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.240000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.480000 ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 46.131199 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 110.055 199.500 124.155 202.460 ;
        RECT 127.955 202.000 128.555 202.300 ;
        RECT 124.555 197.500 135.135 200.460 ;
        RECT 135.555 196.000 143.655 198.960 ;
        RECT 119.055 192.500 124.155 195.460 ;
        RECT 144.055 194.000 150.395 196.960 ;
        RECT 119.905 191.760 121.355 192.500 ;
        RECT 119.505 188.800 123.725 191.760 ;
        RECT 122.705 185.150 125.665 188.750 ;
        RECT 122.705 181.950 129.115 185.050 ;
        RECT 129.405 184.930 132.505 185.480 ;
        RECT 132.955 184.930 136.055 185.310 ;
        RECT 136.535 184.930 139.635 185.340 ;
        RECT 140.115 184.930 143.215 185.470 ;
        RECT 143.695 184.930 146.795 185.450 ;
        RECT 147.275 184.930 150.375 185.440 ;
        RECT 129.405 181.860 150.375 184.930 ;
        RECT 129.405 181.400 132.505 181.860 ;
        RECT 132.955 180.350 136.055 181.860 ;
        RECT 136.535 179.140 139.635 181.860 ;
        RECT 140.115 177.510 143.215 181.860 ;
        RECT 143.695 175.010 146.795 181.860 ;
        RECT 147.275 171.480 150.375 181.860 ;
      LAYER li1 ;
        RECT 111.255 202.280 113.055 202.300 ;
        RECT 110.235 202.110 123.975 202.280 ;
        RECT 110.235 199.850 110.405 202.110 ;
        RECT 111.255 202.100 113.055 202.110 ;
        RECT 111.085 201.540 123.125 201.710 ;
        RECT 110.745 200.480 110.915 201.480 ;
        RECT 123.295 200.480 123.465 201.480 ;
        RECT 111.085 200.250 123.125 200.420 ;
        RECT 123.805 199.850 123.975 202.110 ;
        RECT 125.855 200.280 127.655 200.300 ;
        RECT 110.235 199.680 123.975 199.850 ;
        RECT 124.735 200.110 134.955 200.280 ;
        RECT 124.735 197.850 124.905 200.110 ;
        RECT 125.855 200.100 127.655 200.110 ;
        RECT 125.585 199.540 134.105 199.710 ;
        RECT 125.245 198.480 125.415 199.480 ;
        RECT 134.275 198.480 134.445 199.480 ;
        RECT 125.585 198.250 134.105 198.420 ;
        RECT 134.785 197.850 134.955 200.110 ;
        RECT 136.855 198.780 138.755 198.800 ;
        RECT 124.735 197.680 134.955 197.850 ;
        RECT 135.735 198.610 143.475 198.780 ;
        RECT 135.735 196.350 135.905 198.610 ;
        RECT 136.855 198.600 138.755 198.610 ;
        RECT 136.585 198.040 142.625 198.210 ;
        RECT 136.245 196.980 136.415 197.980 ;
        RECT 142.795 196.980 142.965 197.980 ;
        RECT 136.585 196.750 142.625 196.920 ;
        RECT 143.305 196.350 143.475 198.610 ;
        RECT 145.055 196.780 146.855 196.800 ;
        RECT 135.735 196.180 143.475 196.350 ;
        RECT 144.235 196.610 150.215 196.780 ;
        RECT 119.235 195.110 123.975 195.280 ;
        RECT 119.235 192.850 119.405 195.110 ;
        RECT 120.085 194.540 123.125 194.710 ;
        RECT 119.745 193.480 119.915 194.480 ;
        RECT 123.295 193.480 123.465 194.480 ;
        RECT 120.085 193.250 123.125 193.420 ;
        RECT 123.805 192.850 123.975 195.110 ;
        RECT 144.235 194.350 144.405 196.610 ;
        RECT 145.055 196.600 146.855 196.610 ;
        RECT 145.085 196.040 149.365 196.210 ;
        RECT 144.745 194.980 144.915 195.980 ;
        RECT 149.535 194.980 149.705 195.980 ;
        RECT 145.085 194.750 149.365 194.920 ;
        RECT 150.045 194.350 150.215 196.610 ;
        RECT 144.235 194.180 150.215 194.350 ;
        RECT 119.235 192.680 123.975 192.850 ;
        RECT 119.755 192.650 121.305 192.680 ;
        RECT 120.155 191.580 121.305 191.600 ;
        RECT 119.685 191.410 123.545 191.580 ;
        RECT 119.685 189.150 119.855 191.410 ;
        RECT 120.155 191.400 121.305 191.410 ;
        RECT 120.535 190.840 122.695 191.010 ;
        RECT 120.195 189.780 120.365 190.780 ;
        RECT 122.865 189.780 123.035 190.780 ;
        RECT 120.535 189.550 122.695 189.720 ;
        RECT 123.375 189.150 123.545 191.410 ;
        RECT 119.685 188.980 123.545 189.150 ;
        RECT 123.905 188.570 124.955 188.600 ;
        RECT 122.885 188.400 125.485 188.570 ;
        RECT 122.885 185.500 123.055 188.400 ;
        RECT 123.685 187.890 124.685 188.060 ;
        RECT 123.455 186.180 123.625 187.720 ;
        RECT 124.745 186.180 124.915 187.720 ;
        RECT 123.685 185.840 124.685 186.010 ;
        RECT 125.315 185.500 125.485 188.400 ;
        RECT 122.885 185.330 125.485 185.500 ;
        RECT 123.405 185.300 124.955 185.330 ;
        RECT 129.585 185.130 132.325 185.300 ;
        RECT 123.405 184.870 124.955 184.900 ;
        RECT 127.355 184.870 128.455 184.950 ;
        RECT 122.885 184.700 125.485 184.870 ;
        RECT 122.885 182.300 123.055 184.700 ;
        RECT 123.685 184.190 124.685 184.360 ;
        RECT 123.455 182.980 123.625 184.020 ;
        RECT 124.745 182.980 124.915 184.020 ;
        RECT 123.685 182.640 124.685 182.810 ;
        RECT 125.315 182.300 125.485 184.700 ;
        RECT 122.885 182.130 125.485 182.300 ;
        RECT 125.835 184.700 128.935 184.870 ;
        RECT 129.585 184.850 129.755 185.130 ;
        RECT 129.955 185.050 130.405 185.130 ;
        RECT 125.835 182.300 126.005 184.700 ;
        RECT 126.635 184.190 128.135 184.360 ;
        RECT 126.405 182.980 126.575 184.020 ;
        RECT 128.195 182.980 128.365 184.020 ;
        RECT 126.635 182.640 128.135 182.810 ;
        RECT 128.765 182.300 128.935 184.700 ;
        RECT 129.505 184.450 129.755 184.850 ;
        RECT 130.435 184.560 131.475 184.730 ;
        RECT 125.835 182.130 128.935 182.300 ;
        RECT 129.585 181.750 129.755 184.450 ;
        RECT 130.095 182.380 130.265 184.500 ;
        RECT 131.645 182.380 131.815 184.500 ;
        RECT 130.435 182.150 131.475 182.320 ;
        RECT 132.155 181.750 132.325 185.130 ;
        RECT 129.585 181.580 132.325 181.750 ;
        RECT 133.135 184.960 135.875 185.130 ;
        RECT 133.135 180.700 133.305 184.960 ;
        RECT 135.705 184.820 135.875 184.960 ;
        RECT 136.715 184.990 139.455 185.160 ;
        RECT 133.985 184.390 135.025 184.560 ;
        RECT 133.645 181.330 133.815 184.330 ;
        RECT 135.195 181.330 135.365 184.330 ;
        RECT 135.705 182.060 135.905 184.820 ;
        RECT 133.985 181.100 135.025 181.270 ;
        RECT 135.705 180.700 135.875 182.060 ;
        RECT 133.135 180.530 135.875 180.700 ;
        RECT 136.715 179.490 136.885 184.990 ;
        RECT 139.285 184.820 139.455 184.990 ;
        RECT 140.295 185.120 143.035 185.290 ;
        RECT 137.565 184.420 138.605 184.590 ;
        RECT 137.225 180.120 137.395 184.360 ;
        RECT 138.775 180.120 138.945 184.360 ;
        RECT 139.285 182.060 139.485 184.820 ;
        RECT 137.565 179.890 138.605 180.060 ;
        RECT 139.285 179.490 139.455 182.060 ;
        RECT 136.715 179.320 139.455 179.490 ;
        RECT 140.295 177.860 140.465 185.120 ;
        RECT 142.865 184.820 143.035 185.120 ;
        RECT 143.875 185.100 146.615 185.270 ;
        RECT 141.145 184.550 142.185 184.720 ;
        RECT 140.805 178.490 140.975 184.490 ;
        RECT 142.355 178.490 142.525 184.490 ;
        RECT 142.865 182.060 143.065 184.820 ;
        RECT 141.145 178.260 142.185 178.430 ;
        RECT 142.865 177.860 143.035 182.060 ;
        RECT 140.295 177.690 143.035 177.860 ;
        RECT 143.875 175.360 144.045 185.100 ;
        RECT 146.445 184.820 146.615 185.100 ;
        RECT 147.455 185.090 150.195 185.260 ;
        RECT 144.725 184.530 145.765 184.700 ;
        RECT 144.385 175.990 144.555 184.470 ;
        RECT 145.935 175.990 146.105 184.470 ;
        RECT 146.445 182.060 146.645 184.820 ;
        RECT 144.725 175.760 145.765 175.930 ;
        RECT 146.445 175.360 146.615 182.060 ;
        RECT 143.875 175.190 146.615 175.360 ;
        RECT 147.455 171.830 147.625 185.090 ;
        RECT 148.305 184.520 149.345 184.690 ;
        RECT 147.965 172.460 148.135 184.460 ;
        RECT 149.515 172.460 149.685 184.460 ;
        RECT 150.025 174.900 150.195 185.090 ;
        RECT 148.305 172.230 149.345 172.400 ;
        RECT 150.005 172.150 150.205 174.900 ;
        RECT 150.025 171.830 150.195 172.150 ;
        RECT 147.455 171.660 150.195 171.830 ;
      LAYER met1 ;
        RECT 111.155 205.000 113.155 205.030 ;
        RECT 108.055 203.000 113.155 205.000 ;
        RECT 154.045 204.000 156.445 204.030 ;
        RECT 111.155 202.000 113.155 203.000 ;
        RECT 113.455 202.500 156.445 204.000 ;
        RECT 113.455 202.200 133.555 202.500 ;
        RECT 113.455 202.000 125.455 202.200 ;
        RECT 108.055 201.400 109.055 202.000 ;
        RECT 113.455 201.815 123.055 202.000 ;
        RECT 111.165 201.740 123.055 201.815 ;
        RECT 111.105 201.510 123.105 201.740 ;
        RECT 110.715 201.430 110.945 201.460 ;
        RECT 108.040 201.000 109.055 201.400 ;
        RECT 108.040 200.550 108.950 201.000 ;
        RECT 110.090 200.520 110.945 201.430 ;
        RECT 110.715 200.500 110.945 200.520 ;
        RECT 123.265 201.430 123.495 201.460 ;
        RECT 123.265 200.520 124.140 201.430 ;
        RECT 123.265 200.500 123.495 200.520 ;
        RECT 111.105 200.220 123.105 200.450 ;
        RECT 108.055 199.000 109.055 200.000 ;
        RECT 108.055 198.530 108.895 199.000 ;
        RECT 111.165 198.500 123.045 200.220 ;
        RECT 125.725 200.000 127.785 202.000 ;
        RECT 128.155 201.500 133.555 202.200 ;
        RECT 134.555 201.570 156.445 202.500 ;
        RECT 134.555 201.500 155.555 201.570 ;
        RECT 128.155 201.000 155.555 201.500 ;
        RECT 128.155 200.400 136.455 201.000 ;
        RECT 128.155 199.800 134.015 200.400 ;
        RECT 125.665 199.740 134.015 199.800 ;
        RECT 125.605 199.510 134.085 199.740 ;
        RECT 125.215 199.430 125.445 199.460 ;
        RECT 134.245 199.430 134.475 199.460 ;
        RECT 124.585 198.530 125.445 199.430 ;
        RECT 134.215 198.530 135.055 199.430 ;
        RECT 125.215 198.500 125.445 198.530 ;
        RECT 134.245 198.500 134.475 198.530 ;
        RECT 136.725 198.500 138.785 200.500 ;
        RECT 139.055 200.000 142.055 201.000 ;
        RECT 108.055 197.000 109.055 198.000 ;
        RECT 111.055 197.520 123.045 198.500 ;
        RECT 125.605 198.220 134.085 198.450 ;
        RECT 139.055 198.300 142.515 200.000 ;
        RECT 143.055 199.100 155.555 201.000 ;
        RECT 147.255 198.790 149.255 199.100 ;
        RECT 136.685 198.240 142.515 198.300 ;
        RECT 108.000 196.000 108.870 196.315 ;
        RECT 108.000 195.505 109.055 196.000 ;
        RECT 108.055 195.000 109.055 195.505 ;
        RECT 108.050 194.000 108.860 194.350 ;
        RECT 108.050 193.600 109.055 194.000 ;
        RECT 108.055 193.000 109.055 193.600 ;
        RECT 108.055 191.705 109.055 192.000 ;
        RECT 108.030 191.000 109.055 191.705 ;
        RECT 108.030 190.895 108.780 191.000 ;
        RECT 108.055 189.000 109.055 190.000 ;
        RECT 108.130 188.670 108.880 189.000 ;
        RECT 111.055 188.750 114.055 197.520 ;
        RECT 120.115 197.400 123.045 197.520 ;
        RECT 125.665 197.400 134.015 198.220 ;
        RECT 136.605 198.010 142.605 198.240 ;
        RECT 136.215 197.920 136.445 197.960 ;
        RECT 142.765 197.920 142.995 197.960 ;
        RECT 120.115 196.650 134.015 197.400 ;
        RECT 135.665 197.040 136.485 197.920 ;
        RECT 142.765 197.040 143.615 197.920 ;
        RECT 136.215 197.000 136.445 197.040 ;
        RECT 142.765 197.000 142.995 197.040 ;
        RECT 136.605 196.720 142.605 196.950 ;
        RECT 120.115 196.400 133.955 196.650 ;
        RECT 136.685 196.400 142.515 196.720 ;
        RECT 144.925 196.500 146.985 198.500 ;
        RECT 120.115 195.600 142.515 196.400 ;
        RECT 147.255 196.300 149.265 198.790 ;
        RECT 145.185 196.240 149.265 196.300 ;
        RECT 145.105 196.010 149.345 196.240 ;
        RECT 144.715 195.910 144.945 195.960 ;
        RECT 120.115 194.740 123.045 195.600 ;
        RECT 132.155 194.840 142.515 195.600 ;
        RECT 144.110 195.040 144.945 195.910 ;
        RECT 144.715 195.000 144.945 195.040 ;
        RECT 149.505 195.910 149.735 195.960 ;
        RECT 149.505 195.040 150.320 195.910 ;
        RECT 149.505 195.000 149.735 195.040 ;
        RECT 120.105 194.510 123.105 194.740 ;
        RECT 132.155 194.600 142.455 194.840 ;
        RECT 145.105 194.720 149.345 194.950 ;
        RECT 119.715 194.380 119.945 194.460 ;
        RECT 119.180 193.570 119.945 194.380 ;
        RECT 119.715 193.500 119.945 193.570 ;
        RECT 123.265 194.380 123.495 194.460 ;
        RECT 123.265 193.570 124.080 194.380 ;
        RECT 137.675 194.190 141.935 194.600 ;
        RECT 145.185 194.190 149.265 194.720 ;
        RECT 123.265 193.500 123.495 193.570 ;
        RECT 120.105 193.220 123.105 193.450 ;
        RECT 121.555 193.050 123.055 193.220 ;
        RECT 119.655 191.300 121.405 193.000 ;
        RECT 121.555 191.800 136.705 193.050 ;
        RECT 137.675 192.200 149.265 194.190 ;
        RECT 150.655 191.800 155.555 199.100 ;
        RECT 121.555 191.700 155.555 191.800 ;
        RECT 121.555 191.040 122.605 191.700 ;
        RECT 122.785 191.680 155.555 191.700 ;
        RECT 120.555 190.810 122.675 191.040 ;
        RECT 123.955 190.800 125.055 190.850 ;
        RECT 120.165 190.630 120.395 190.760 ;
        RECT 122.835 190.630 123.065 190.760 ;
        RECT 120.135 190.600 120.780 190.630 ;
        RECT 120.105 189.955 120.810 190.600 ;
        RECT 120.135 189.925 120.780 189.955 ;
        RECT 122.430 189.925 123.075 190.630 ;
        RECT 120.165 189.800 120.395 189.925 ;
        RECT 122.835 189.800 123.065 189.925 ;
        RECT 120.555 189.520 122.675 189.750 ;
        RECT 123.925 189.700 125.085 190.800 ;
        RECT 120.605 188.750 122.605 189.520 ;
        RECT 108.055 187.000 109.055 188.000 ;
        RECT 111.055 187.600 122.605 188.750 ;
        RECT 123.805 188.350 125.055 189.700 ;
        RECT 123.805 188.090 124.505 188.120 ;
        RECT 123.705 187.860 124.665 188.090 ;
        RECT 123.425 187.600 123.655 187.700 ;
        RECT 108.130 186.520 108.880 187.000 ;
        RECT 111.055 186.750 123.655 187.600 ;
        RECT 123.805 187.480 124.505 187.860 ;
        RECT 124.715 187.600 124.945 187.700 ;
        RECT 128.805 187.600 155.555 191.680 ;
        RECT 108.055 185.000 109.055 186.000 ;
        RECT 108.080 184.670 108.830 185.000 ;
        RECT 108.055 183.625 109.055 184.000 ;
        RECT 108.050 183.000 109.055 183.625 ;
        RECT 108.050 182.875 108.860 183.000 ;
        RECT 108.055 181.000 109.055 182.000 ;
        RECT 108.080 180.795 108.830 181.000 ;
        RECT 108.055 179.625 109.055 180.000 ;
        RECT 108.000 179.000 109.055 179.625 ;
        RECT 108.000 178.875 108.810 179.000 ;
        RECT 108.055 177.760 109.055 178.000 ;
        RECT 108.030 177.000 109.055 177.760 ;
        RECT 108.030 176.950 108.780 177.000 ;
        RECT 108.055 175.000 109.055 176.000 ;
        RECT 108.100 174.825 108.910 175.000 ;
        RECT 108.055 173.825 109.055 174.000 ;
        RECT 108.000 173.075 109.055 173.825 ;
        RECT 108.055 173.000 109.055 173.075 ;
        RECT 111.055 172.000 114.055 186.750 ;
        RECT 120.605 186.300 123.655 186.750 ;
        RECT 123.835 186.370 124.475 187.480 ;
        RECT 120.605 183.900 122.605 186.300 ;
        RECT 123.425 186.200 123.655 186.300 ;
        RECT 123.805 186.040 124.505 186.370 ;
        RECT 124.715 186.310 155.555 187.600 ;
        RECT 124.715 186.300 150.575 186.310 ;
        RECT 124.715 186.200 124.945 186.300 ;
        RECT 123.705 185.810 124.665 186.040 ;
        RECT 123.805 185.730 124.505 185.810 ;
        RECT 123.305 184.650 125.055 185.550 ;
        RECT 123.850 184.390 124.565 184.425 ;
        RECT 123.705 184.160 124.665 184.390 ;
        RECT 123.425 183.900 123.655 184.000 ;
        RECT 120.605 183.100 123.655 183.900 ;
        RECT 123.850 183.770 124.565 184.160 ;
        RECT 124.715 183.900 124.945 184.000 ;
        RECT 125.255 183.900 126.030 186.300 ;
        RECT 127.325 186.000 128.485 186.150 ;
        RECT 127.325 185.100 130.505 186.000 ;
        RECT 127.305 185.000 130.505 185.100 ;
        RECT 127.305 184.650 128.505 185.000 ;
        RECT 127.230 184.390 127.980 184.405 ;
        RECT 129.405 184.400 129.855 185.000 ;
        RECT 130.655 184.760 131.455 186.300 ;
        RECT 132.155 184.920 133.305 184.930 ;
        RECT 132.115 184.910 133.355 184.920 ;
        RECT 126.655 184.160 128.115 184.390 ;
        RECT 130.065 184.225 130.295 184.480 ;
        RECT 130.455 184.450 131.455 184.760 ;
        RECT 131.615 184.255 131.845 184.480 ;
        RECT 126.375 183.900 126.605 184.000 ;
        RECT 123.425 183.000 123.655 183.100 ;
        RECT 123.850 182.840 124.565 183.230 ;
        RECT 124.715 183.050 126.755 183.900 ;
        RECT 127.230 183.595 127.980 184.160 ;
        RECT 124.715 183.000 124.945 183.050 ;
        RECT 126.375 183.000 126.605 183.050 ;
        RECT 126.950 182.840 127.760 183.225 ;
        RECT 128.165 183.000 129.305 184.000 ;
        RECT 129.500 183.475 130.310 184.225 ;
        RECT 128.255 182.950 129.305 183.000 ;
        RECT 123.705 182.610 124.665 182.840 ;
        RECT 126.655 182.610 128.115 182.840 ;
        RECT 123.850 182.575 124.565 182.610 ;
        RECT 126.950 182.475 127.760 182.610 ;
        RECT 128.405 181.210 129.305 182.950 ;
        RECT 129.530 182.395 130.310 183.475 ;
        RECT 131.130 182.500 131.865 184.255 ;
        RECT 131.615 182.400 131.845 182.500 ;
        RECT 128.395 172.000 129.395 181.210 ;
        RECT 130.455 172.000 131.455 182.350 ;
        RECT 132.085 181.860 133.355 184.910 ;
        RECT 133.975 184.390 135.015 186.300 ;
        RECT 136.255 186.280 138.585 186.300 ;
        RECT 135.735 184.920 136.885 184.930 ;
        RECT 135.695 184.910 136.935 184.920 ;
        RECT 134.005 184.360 135.005 184.390 ;
        RECT 133.615 184.105 133.845 184.310 ;
        RECT 135.165 184.135 135.395 184.310 ;
        RECT 133.540 183.355 134.350 184.105 ;
        RECT 133.615 181.350 133.845 183.355 ;
        RECT 134.670 183.325 135.420 184.135 ;
        RECT 135.165 181.350 135.395 183.325 ;
        RECT 135.665 181.860 136.935 184.910 ;
        RECT 137.585 184.390 138.585 186.280 ;
        RECT 139.315 184.920 140.465 184.930 ;
        RECT 139.275 184.910 140.515 184.920 ;
        RECT 137.195 184.165 137.425 184.340 ;
        RECT 138.745 184.195 138.975 184.340 ;
        RECT 137.145 183.415 137.955 184.165 ;
        RECT 134.005 181.250 135.005 181.300 ;
        RECT 134.005 172.000 135.015 181.250 ;
        RECT 137.195 181.065 137.425 183.415 ;
        RECT 138.280 183.385 139.030 184.195 ;
        RECT 137.150 180.315 137.960 181.065 ;
        RECT 138.745 180.985 138.975 183.385 ;
        RECT 139.245 181.860 140.515 184.910 ;
        RECT 141.155 184.750 142.155 186.300 ;
        RECT 142.895 184.920 144.045 184.930 ;
        RECT 142.855 184.910 144.095 184.920 ;
        RECT 141.155 184.550 142.165 184.750 ;
        RECT 141.165 184.520 142.165 184.550 ;
        RECT 140.775 184.295 141.005 184.470 ;
        RECT 142.325 184.325 142.555 184.470 ;
        RECT 140.705 183.545 141.515 184.295 ;
        RECT 137.195 180.140 137.425 180.315 ;
        RECT 138.250 180.235 139.060 180.985 ;
        RECT 138.745 180.140 138.975 180.235 ;
        RECT 137.585 179.860 138.585 180.090 ;
        RECT 137.595 172.000 138.525 179.860 ;
        RECT 140.775 179.455 141.005 183.545 ;
        RECT 141.860 183.515 142.610 184.325 ;
        RECT 140.740 178.645 141.490 179.455 ;
        RECT 142.325 179.425 142.555 183.515 ;
        RECT 142.825 181.860 144.095 184.910 ;
        RECT 144.755 184.730 145.755 186.300 ;
        RECT 146.475 184.920 147.625 184.930 ;
        RECT 146.435 184.910 147.675 184.920 ;
        RECT 144.745 184.540 145.755 184.730 ;
        RECT 144.745 184.500 145.745 184.540 ;
        RECT 144.355 184.315 144.585 184.450 ;
        RECT 145.905 184.345 146.135 184.450 ;
        RECT 144.265 183.565 145.075 184.315 ;
        RECT 141.830 178.675 142.640 179.425 ;
        RECT 140.775 178.510 141.005 178.645 ;
        RECT 142.325 178.510 142.555 178.675 ;
        RECT 141.175 178.460 142.105 178.480 ;
        RECT 141.165 178.230 142.165 178.460 ;
        RECT 141.175 172.000 142.105 178.230 ;
        RECT 144.355 176.925 144.585 183.565 ;
        RECT 145.430 183.535 146.180 184.345 ;
        RECT 144.310 176.115 145.060 176.925 ;
        RECT 145.905 176.895 146.135 183.535 ;
        RECT 146.405 181.860 147.675 184.910 ;
        RECT 148.315 184.720 149.315 186.300 ;
        RECT 148.315 184.510 149.325 184.720 ;
        RECT 148.325 184.490 149.325 184.510 ;
        RECT 147.935 184.285 148.165 184.440 ;
        RECT 149.485 184.315 149.715 184.440 ;
        RECT 147.865 183.535 148.675 184.285 ;
        RECT 145.400 176.145 146.210 176.895 ;
        RECT 144.355 176.010 144.585 176.115 ;
        RECT 145.905 176.010 146.135 176.145 ;
        RECT 144.745 175.730 145.745 175.960 ;
        RECT 144.755 172.000 145.685 175.730 ;
        RECT 147.935 173.405 148.165 183.535 ;
        RECT 149.030 183.505 149.780 184.315 ;
        RECT 147.900 172.595 148.650 173.405 ;
        RECT 149.485 173.375 149.715 183.505 ;
        RECT 149.000 172.625 149.810 173.375 ;
        RECT 147.935 172.480 148.165 172.595 ;
        RECT 149.485 172.480 149.715 172.625 ;
        RECT 148.325 172.200 149.325 172.430 ;
        RECT 104.270 171.280 147.055 172.000 ;
        RECT 148.335 171.280 149.315 172.200 ;
        RECT 149.955 171.850 151.605 175.000 ;
        RECT 150.205 171.700 151.605 171.850 ;
        RECT 104.270 170.260 149.315 171.280 ;
        RECT 104.270 169.000 147.055 170.260 ;
      LAYER met2 ;
        RECT 104.800 204.770 152.765 205.000 ;
        RECT 104.775 204.750 152.765 204.770 ;
        RECT 104.750 203.250 152.765 204.750 ;
        RECT 104.775 203.230 152.765 203.250 ;
        RECT 104.800 203.000 152.765 203.230 ;
        RECT 105.755 201.400 109.065 202.170 ;
        RECT 105.755 200.975 124.610 201.400 ;
        RECT 108.070 200.550 124.610 200.975 ;
        RECT 108.070 200.520 108.920 200.550 ;
        RECT 105.755 199.400 109.075 200.170 ;
        RECT 125.755 199.970 127.755 203.000 ;
        RECT 105.755 198.975 135.090 199.400 ;
        RECT 108.025 198.560 135.090 198.975 ;
        RECT 136.755 198.470 138.755 203.000 ;
        RECT 105.755 197.890 109.035 198.170 ;
        RECT 105.755 197.070 143.735 197.890 ;
        RECT 105.755 196.975 109.035 197.070 ;
        RECT 144.955 196.470 146.955 203.000 ;
        RECT 108.030 196.315 108.840 196.345 ;
        RECT 108.030 196.170 126.040 196.315 ;
        RECT 105.755 195.880 126.040 196.170 ;
        RECT 105.755 195.505 150.480 195.880 ;
        RECT 105.755 194.975 109.075 195.505 ;
        RECT 125.230 195.070 150.480 195.505 ;
        RECT 108.080 194.350 108.830 194.380 ;
        RECT 108.080 194.170 124.110 194.350 ;
        RECT 105.755 193.600 124.110 194.170 ;
        RECT 105.755 192.975 109.065 193.600 ;
        RECT 150.765 192.850 152.765 203.000 ;
        RECT 153.900 201.600 157.300 204.000 ;
        RECT 105.755 191.675 109.095 192.170 ;
        RECT 105.755 190.975 110.780 191.675 ;
        RECT 119.775 191.450 152.765 192.850 ;
        RECT 108.000 190.925 110.780 190.975 ;
        RECT 110.030 190.650 110.780 190.925 ;
        RECT 105.755 189.450 109.105 190.170 ;
        RECT 110.030 189.900 123.230 190.650 ;
        RECT 123.955 189.670 125.055 191.450 ;
        RECT 105.755 188.975 124.480 189.450 ;
        RECT 108.055 188.700 124.480 188.975 ;
        RECT 105.755 187.300 109.095 188.170 ;
        RECT 105.755 186.975 120.430 187.300 ;
        RECT 108.055 186.550 120.430 186.975 ;
        RECT 105.755 185.450 109.075 186.170 ;
        RECT 105.755 184.975 118.930 185.450 ;
        RECT 108.050 184.700 118.930 184.975 ;
        RECT 105.755 183.075 109.075 184.170 ;
        RECT 105.755 182.975 117.380 183.075 ;
        RECT 108.055 182.325 117.380 182.975 ;
        RECT 105.755 181.575 109.085 182.170 ;
        RECT 105.755 180.975 115.680 181.575 ;
        RECT 108.050 180.825 115.680 180.975 ;
        RECT 114.930 180.250 115.680 180.825 ;
        RECT 116.630 181.225 117.380 182.325 ;
        RECT 118.180 182.275 118.930 184.700 ;
        RECT 119.680 185.175 120.430 186.550 ;
        RECT 123.835 185.700 124.475 188.700 ;
        RECT 127.355 187.680 128.455 191.450 ;
        RECT 150.755 187.680 152.765 191.450 ;
        RECT 127.355 186.280 152.765 187.680 ;
        RECT 119.680 184.425 124.580 185.175 ;
        RECT 127.355 185.020 128.455 186.280 ;
        RECT 119.680 184.400 120.430 184.425 ;
        RECT 123.880 182.545 124.535 184.425 ;
        RECT 126.780 182.275 128.030 184.375 ;
        RECT 129.530 183.275 131.865 184.325 ;
        RECT 132.355 183.575 133.105 186.280 ;
        RECT 133.555 184.105 135.440 184.245 ;
        RECT 129.500 182.625 131.865 183.275 ;
        RECT 118.180 181.525 128.030 182.275 ;
        RECT 129.530 182.550 131.865 182.625 ;
        RECT 133.555 183.355 135.450 184.105 ;
        RECT 135.935 183.575 136.685 186.280 ;
        RECT 137.175 184.165 137.925 184.245 ;
        RECT 137.175 183.415 139.060 184.165 ;
        RECT 139.515 183.575 140.265 186.280 ;
        RECT 140.735 184.295 141.485 184.325 ;
        RECT 140.735 183.545 142.640 184.295 ;
        RECT 143.095 183.575 143.845 186.280 ;
        RECT 144.295 184.315 145.045 184.345 ;
        RECT 144.295 183.565 146.210 184.315 ;
        RECT 146.675 183.575 147.425 186.280 ;
        RECT 147.895 184.285 148.645 184.315 ;
        RECT 129.530 182.500 131.130 182.550 ;
        RECT 129.530 181.225 130.280 182.500 ;
        RECT 116.630 180.475 130.280 181.225 ;
        RECT 133.555 182.215 134.320 183.355 ;
        RECT 134.690 182.215 135.440 183.355 ;
        RECT 133.555 181.465 135.440 182.215 ;
        RECT 137.175 182.565 137.925 183.415 ;
        RECT 133.555 180.250 134.305 181.465 ;
        RECT 137.175 180.985 137.930 182.565 ;
        RECT 138.280 180.985 139.030 183.415 ;
        RECT 105.755 178.990 109.055 180.170 ;
        RECT 114.930 179.500 134.330 180.250 ;
        RECT 137.175 180.235 139.030 180.985 ;
        RECT 137.175 178.990 137.925 180.235 ;
        RECT 138.280 180.205 139.030 180.235 ;
        RECT 140.735 179.425 141.485 183.545 ;
        RECT 141.860 179.425 142.610 183.545 ;
        RECT 105.755 178.975 137.925 178.990 ;
        RECT 108.030 178.240 137.925 178.975 ;
        RECT 140.710 178.675 142.610 179.425 ;
        RECT 105.745 177.730 109.075 177.970 ;
        RECT 140.735 177.730 141.485 178.675 ;
        RECT 141.860 178.645 142.610 178.675 ;
        RECT 105.745 176.980 141.485 177.730 ;
        RECT 105.745 176.775 109.075 176.980 ;
        RECT 144.295 176.895 145.045 183.565 ;
        RECT 145.430 176.895 146.180 183.565 ;
        RECT 105.755 175.150 109.085 176.170 ;
        RECT 144.280 176.145 146.180 176.895 ;
        RECT 144.295 175.150 145.045 176.145 ;
        RECT 145.430 176.115 146.180 176.145 ;
        RECT 147.895 183.535 149.810 184.285 ;
        RECT 105.755 174.975 145.045 175.150 ;
        RECT 108.130 174.400 145.045 174.975 ;
        RECT 105.755 172.975 109.075 174.170 ;
        RECT 147.895 173.375 148.645 183.535 ;
        RECT 149.030 173.375 149.780 183.535 ;
        RECT 150.765 173.550 152.765 186.280 ;
        RECT 108.030 172.125 108.780 172.975 ;
        RECT 147.870 172.625 149.780 173.375 ;
        RECT 147.895 172.125 148.645 172.625 ;
        RECT 149.030 172.595 149.780 172.625 ;
        RECT 150.175 172.150 152.765 173.550 ;
        RECT 104.300 172.000 107.300 172.030 ;
        RECT 102.600 169.000 107.300 172.000 ;
        RECT 108.030 171.375 148.645 172.125 ;
        RECT 150.765 172.100 152.765 172.150 ;
        RECT 147.895 171.290 148.645 171.375 ;
        RECT 104.300 168.970 107.300 169.000 ;
      LAYER met3 ;
        RECT 87.015 204.750 88.505 204.775 ;
        RECT 87.010 203.250 106.250 204.750 ;
        RECT 156.425 203.280 157.300 203.305 ;
        RECT 87.015 203.225 88.505 203.250 ;
        RECT 156.420 202.395 157.305 203.280 ;
        RECT 156.425 202.370 157.300 202.395 ;
        RECT 105.380 201.140 106.780 202.000 ;
        RECT 105.380 199.140 106.780 200.000 ;
        RECT 105.380 197.140 106.780 198.000 ;
        RECT 105.380 195.140 106.780 196.000 ;
        RECT 105.380 193.140 106.780 194.000 ;
        RECT 105.380 191.140 106.780 192.000 ;
        RECT 105.380 189.140 106.780 190.000 ;
        RECT 105.380 187.140 106.780 188.000 ;
        RECT 105.380 185.140 106.780 186.000 ;
        RECT 105.380 183.140 106.780 184.000 ;
        RECT 105.380 181.140 106.780 182.000 ;
        RECT 105.380 179.140 106.780 180.000 ;
        RECT 105.370 176.940 106.770 177.800 ;
        RECT 105.380 175.140 106.780 176.000 ;
        RECT 105.380 173.140 106.780 174.000 ;
        RECT 44.755 171.250 46.245 171.275 ;
        RECT 44.750 169.750 104.250 171.250 ;
        RECT 44.755 169.725 46.245 169.750 ;
      LAYER met4 ;
        RECT 3.990 223.540 4.290 224.760 ;
        RECT 7.670 223.540 7.970 224.760 ;
        RECT 11.350 223.540 11.650 224.760 ;
        RECT 15.030 223.540 15.330 224.760 ;
        RECT 18.710 223.540 19.010 224.760 ;
        RECT 22.390 223.540 22.690 224.760 ;
        RECT 26.070 223.540 26.370 224.760 ;
        RECT 29.750 223.540 30.050 224.760 ;
        RECT 33.430 223.540 33.730 224.760 ;
        RECT 37.110 223.540 37.410 224.760 ;
        RECT 40.790 223.540 41.090 224.760 ;
        RECT 44.470 223.540 44.770 224.760 ;
        RECT 48.150 223.540 48.450 224.760 ;
        RECT 51.830 223.540 52.130 224.760 ;
        RECT 55.510 223.540 55.810 224.760 ;
        RECT 59.190 223.540 59.490 224.760 ;
        RECT 62.870 223.540 63.170 224.760 ;
        RECT 66.550 223.540 66.850 224.760 ;
        RECT 70.230 223.540 70.530 224.760 ;
        RECT 73.910 223.540 74.210 224.760 ;
        RECT 77.590 223.540 77.890 224.760 ;
        RECT 81.270 223.540 81.570 224.760 ;
        RECT 84.950 223.540 85.250 224.760 ;
        RECT 88.630 223.540 88.930 224.760 ;
        RECT 3.990 223.240 88.930 223.540 ;
        RECT 29.750 220.420 30.050 223.240 ;
        RECT 49.550 220.760 49.850 223.240 ;
        RECT 51.830 223.210 52.130 223.240 ;
        RECT 29.750 220.120 49.000 220.420 ;
        RECT 50.500 203.250 88.510 204.750 ;
        RECT 92.310 173.720 92.610 224.760 ;
        RECT 95.990 218.720 96.290 224.760 ;
        RECT 92.990 218.600 96.290 218.720 ;
        RECT 92.990 218.420 96.280 218.600 ;
        RECT 92.990 175.720 93.290 218.420 ;
        RECT 99.670 218.020 99.970 224.760 ;
        RECT 93.690 217.720 99.980 218.020 ;
        RECT 93.690 177.530 93.990 217.720 ;
        RECT 99.670 217.710 99.970 217.720 ;
        RECT 103.350 217.320 103.650 224.760 ;
        RECT 94.410 217.020 103.650 217.320 ;
        RECT 94.410 179.710 94.710 217.020 ;
        RECT 103.350 217.010 103.650 217.020 ;
        RECT 107.030 216.660 107.330 224.760 ;
        RECT 95.230 216.360 107.330 216.660 ;
        RECT 95.230 181.710 95.530 216.360 ;
        RECT 110.710 216.050 111.010 224.760 ;
        RECT 96.030 215.750 111.010 216.050 ;
        RECT 96.030 183.710 96.330 215.750 ;
        RECT 114.390 215.400 114.690 224.760 ;
        RECT 96.710 215.100 114.690 215.400 ;
        RECT 96.710 185.700 97.010 215.100 ;
        RECT 118.070 214.780 118.370 224.760 ;
        RECT 115.070 214.590 118.370 214.780 ;
        RECT 97.440 214.290 118.370 214.590 ;
        RECT 97.440 187.690 97.740 214.290 ;
        RECT 121.750 213.960 122.050 224.760 ;
        RECT 98.140 213.660 122.050 213.960 ;
        RECT 98.140 189.700 98.440 213.660 ;
        RECT 125.430 213.150 125.730 224.760 ;
        RECT 98.910 212.850 125.730 213.150 ;
        RECT 98.910 191.750 99.210 212.850 ;
        RECT 129.110 212.190 129.410 224.760 ;
        RECT 99.600 211.890 129.410 212.190 ;
        RECT 99.600 193.710 99.900 211.890 ;
        RECT 132.790 211.330 133.090 224.760 ;
        RECT 100.240 211.030 133.090 211.330 ;
        RECT 100.240 195.710 100.540 211.030 ;
        RECT 136.470 210.480 136.770 224.760 ;
        RECT 100.930 210.180 136.770 210.480 ;
        RECT 100.930 197.720 101.230 210.180 ;
        RECT 140.150 209.790 140.450 224.760 ;
        RECT 101.680 209.490 140.450 209.790 ;
        RECT 101.680 199.720 101.980 209.490 ;
        RECT 143.830 209.040 144.130 224.760 ;
        RECT 102.370 208.740 144.130 209.040 ;
        RECT 102.370 201.670 102.670 208.740 ;
        RECT 147.510 208.210 147.810 224.760 ;
        RECT 103.090 207.910 147.810 208.210 ;
        RECT 103.090 206.560 103.390 207.910 ;
        RECT 105.645 201.720 105.975 201.735 ;
        RECT 104.920 201.670 105.975 201.720 ;
        RECT 102.370 201.420 105.975 201.670 ;
        RECT 102.370 201.370 105.180 201.420 ;
        RECT 105.645 201.405 105.975 201.420 ;
        RECT 105.645 199.720 105.975 199.735 ;
        RECT 101.680 199.420 105.975 199.720 ;
        RECT 105.645 199.405 105.975 199.420 ;
        RECT 105.645 197.720 105.975 197.735 ;
        RECT 100.930 197.420 105.975 197.720 ;
        RECT 105.645 197.405 105.975 197.420 ;
        RECT 105.645 195.720 105.975 195.735 ;
        RECT 104.920 195.710 105.975 195.720 ;
        RECT 100.240 195.420 105.975 195.710 ;
        RECT 100.240 195.410 105.260 195.420 ;
        RECT 105.645 195.405 105.975 195.420 ;
        RECT 105.645 193.720 105.975 193.735 ;
        RECT 104.920 193.710 105.975 193.720 ;
        RECT 99.600 193.420 105.975 193.710 ;
        RECT 99.600 193.410 105.240 193.420 ;
        RECT 105.645 193.405 105.975 193.420 ;
        RECT 98.910 191.720 105.180 191.750 ;
        RECT 105.645 191.720 105.975 191.735 ;
        RECT 98.910 191.450 105.975 191.720 ;
        RECT 104.920 191.420 105.975 191.450 ;
        RECT 105.645 191.405 105.975 191.420 ;
        RECT 105.645 189.720 105.975 189.735 ;
        RECT 104.920 189.700 105.975 189.720 ;
        RECT 98.140 189.420 105.975 189.700 ;
        RECT 98.140 189.400 105.260 189.420 ;
        RECT 105.645 189.405 105.975 189.420 ;
        RECT 105.645 187.720 105.975 187.735 ;
        RECT 104.920 187.690 105.975 187.720 ;
        RECT 97.440 187.420 105.975 187.690 ;
        RECT 97.440 187.390 105.130 187.420 ;
        RECT 105.645 187.405 105.975 187.420 ;
        RECT 105.645 185.720 105.975 185.735 ;
        RECT 104.920 185.700 105.975 185.720 ;
        RECT 96.710 185.420 105.975 185.700 ;
        RECT 96.710 185.400 105.180 185.420 ;
        RECT 105.645 185.405 105.975 185.420 ;
        RECT 105.645 183.720 105.975 183.735 ;
        RECT 104.920 183.710 105.975 183.720 ;
        RECT 96.030 183.420 105.975 183.710 ;
        RECT 96.030 183.410 105.190 183.420 ;
        RECT 105.645 183.405 105.975 183.420 ;
        RECT 105.645 181.720 105.975 181.735 ;
        RECT 104.920 181.710 105.975 181.720 ;
        RECT 95.230 181.420 105.975 181.710 ;
        RECT 95.230 181.410 105.210 181.420 ;
        RECT 105.645 181.405 105.975 181.420 ;
        RECT 105.645 179.720 105.975 179.735 ;
        RECT 104.920 179.710 105.975 179.720 ;
        RECT 94.410 179.420 105.975 179.710 ;
        RECT 94.410 179.410 105.180 179.420 ;
        RECT 105.645 179.405 105.975 179.420 ;
        RECT 93.690 177.520 105.300 177.530 ;
        RECT 105.635 177.520 105.965 177.535 ;
        RECT 93.690 177.230 105.965 177.520 ;
        RECT 104.910 177.220 105.965 177.230 ;
        RECT 105.635 177.205 105.965 177.220 ;
        RECT 105.645 175.720 105.975 175.735 ;
        RECT 92.990 175.420 105.975 175.720 ;
        RECT 92.990 175.390 93.290 175.420 ;
        RECT 105.645 175.405 105.975 175.420 ;
        RECT 105.645 173.720 105.975 173.735 ;
        RECT 92.310 173.420 105.975 173.720 ;
        RECT 105.645 173.405 105.975 173.420 ;
        RECT 2.500 169.750 46.250 171.250 ;
        RECT 156.420 1.000 157.305 203.280 ;
  END
END tt_um_rejunity_analog_dac_ay8913
END LIBRARY

