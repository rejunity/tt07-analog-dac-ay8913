magic
tech sky130A
timestamp 1716300029
<< pwell >>
rect -310 -155 310 155
<< nmoslvt >>
rect -212 -50 212 50
<< ndiff >>
rect -241 44 -212 50
rect -241 -44 -235 44
rect -218 -44 -212 44
rect -241 -50 -212 -44
rect 212 44 241 50
rect 212 -44 218 44
rect 235 -44 241 44
rect 212 -50 241 -44
<< ndiffc >>
rect -235 -44 -218 44
rect 218 -44 235 44
<< psubdiff >>
rect -292 120 -244 137
rect 244 120 292 137
rect -292 89 -275 120
rect 275 89 292 120
rect -292 -120 -275 -89
rect 275 -120 292 -89
rect -292 -137 -244 -120
rect 244 -137 292 -120
<< psubdiffcont >>
rect -244 120 244 137
rect -292 -89 -275 89
rect 275 -89 292 89
rect -244 -137 244 -120
<< poly >>
rect -212 86 212 94
rect -212 69 -204 86
rect 204 69 212 86
rect -212 50 212 69
rect -212 -69 212 -50
rect -212 -86 -204 -69
rect 204 -86 212 -69
rect -212 -94 212 -86
<< polycont >>
rect -204 69 204 86
rect -204 -86 204 -69
<< locali >>
rect -292 120 -244 137
rect 244 120 292 137
rect -292 89 -275 120
rect 275 89 292 120
rect -212 69 -204 86
rect 204 69 212 86
rect -235 44 -218 52
rect -235 -52 -218 -44
rect 218 44 235 52
rect 218 -52 235 -44
rect -212 -86 -204 -69
rect 204 -86 212 -69
rect -292 -120 -275 -89
rect 275 -120 292 -89
rect -292 -137 -244 -120
rect 244 -137 292 -120
<< viali >>
rect -204 69 204 86
rect -235 -44 -218 44
rect 218 -44 235 44
rect -204 -86 204 -69
<< metal1 >>
rect -210 86 210 89
rect -210 69 -204 86
rect 204 69 210 86
rect -210 66 210 69
rect -238 44 -215 50
rect -238 -44 -235 44
rect -218 -44 -215 44
rect -238 -50 -215 -44
rect 215 44 238 50
rect 215 -44 218 44
rect 235 -44 238 44
rect 215 -50 238 -44
rect -210 -69 210 -66
rect -210 -86 -204 -69
rect 204 -86 210 -69
rect -210 -89 210 -86
<< properties >>
string FIXED_BBOX -283 -128 283 128
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1.0 l 4.24 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
