** sch_path: /Users/rej/Dev/TinyTapeout/tt07-analog-dac-ay8193.git/xschem/dac_16nfet.sch
.subckt dac_16nfet VDD AT0 AT1 AT2 AT3 AT4 AT5 AT6 AT7 AT8 AT9 AT10 AT11 AT12 AT13 AT14 OUT VSS
*.PININFO AT12:I AT13:I VDD:B VSS:B OUT:O AT14:I AT4:I AT5:I AT6:I AT7:I AT8:I AT9:I AT10:I AT11:I AT0:I AT1:I AT2:I AT3:I
XM4 VDD AT0 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=12 nf=1 m=1
XM14 VDD AT1 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=8.484 nf=1 m=1
XM15 VDD AT2 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=6 nf=1 m=1
XM16 VDD AT3 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=4.24 nf=1 m=1
XM9 VDD AT4 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM10 VDD AT5 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=2.12 nf=1 m=1
XM12 VDD AT7 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XM1 VDD AT14 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=12 W=1 nf=1 m=1
XM2 VDD AT13 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=8.484 W=1 nf=1 m=1
XM3 VDD AT12 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=6 W=1 nf=1 m=1
XM5 VDD AT11 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=4.24 W=1 nf=1 m=1
XM6 VDD AT10 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=3 W=1 nf=1 m=1
XM7 VDD AT9 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=2.12 W=1 nf=1 m=1
XM8 VDD AT6 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=1.5 nf=1 m=1
XM11 VDD AT8 OUT VSS sky130_fd_pr__nfet_01v8_lvt L=1.5 W=1 nf=1 m=1
.ends
.end
