magic
tech sky130A
timestamp 1716300029
<< pwell >>
rect -148 -529 148 529
<< nmoslvt >>
rect -50 -424 50 424
<< ndiff >>
rect -79 418 -50 424
rect -79 -418 -73 418
rect -56 -418 -50 418
rect -79 -424 -50 -418
rect 50 418 79 424
rect 50 -418 56 418
rect 73 -418 79 418
rect 50 -424 79 -418
<< ndiffc >>
rect -73 -418 -56 418
rect 56 -418 73 418
<< psubdiff >>
rect -130 494 -82 511
rect 82 494 130 511
rect -130 463 -113 494
rect 113 463 130 494
rect -130 -494 -113 -463
rect 113 -494 130 -463
rect -130 -511 -82 -494
rect 82 -511 130 -494
<< psubdiffcont >>
rect -82 494 82 511
rect -130 -463 -113 463
rect 113 -463 130 463
rect -82 -511 82 -494
<< poly >>
rect -50 460 50 468
rect -50 443 -42 460
rect 42 443 50 460
rect -50 424 50 443
rect -50 -443 50 -424
rect -50 -460 -42 -443
rect 42 -460 50 -443
rect -50 -468 50 -460
<< polycont >>
rect -42 443 42 460
rect -42 -460 42 -443
<< locali >>
rect -130 494 -82 511
rect 82 494 130 511
rect -130 463 -113 494
rect 113 463 130 494
rect -50 443 -42 460
rect 42 443 50 460
rect -73 418 -56 426
rect -73 -426 -56 -418
rect 56 418 73 426
rect 56 -426 73 -418
rect -50 -460 -42 -443
rect 42 -460 50 -443
rect -130 -494 -113 -463
rect 113 -494 130 -463
rect -130 -511 -82 -494
rect 82 -511 130 -494
<< viali >>
rect -42 443 42 460
rect -73 -418 -56 418
rect 56 -418 73 418
rect -42 -460 42 -443
<< metal1 >>
rect -48 460 48 463
rect -48 443 -42 460
rect 42 443 48 460
rect -48 440 48 443
rect -76 418 -53 424
rect -76 -418 -73 418
rect -56 -418 -53 418
rect -76 -424 -53 -418
rect 53 418 76 424
rect 53 -418 56 418
rect 73 -418 76 418
rect 53 -424 76 -418
rect -48 -443 48 -440
rect -48 -460 -42 -443
rect 42 -460 48 -443
rect -48 -463 48 -460
<< properties >>
string FIXED_BBOX -121 -502 121 502
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8.484 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
